��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8F�]��M����B��9DI�Z6�`��c���d
Z�T�:u���V_�g�kkA����_��{]����&	�N�L���r�0�5C؜_]W��c���>&w�@Ⴉ:3��^�!At�<l�LwT�*��A�cG��<��Nn���� <V�s	�`�����dWلv����n��]���4�H�"�>'D��������@2�E�WZ\~`� c�n����j�z����C�b�HMǽ��䢞|�z%A�P� �+M��0�9�'�IP}ad2��)��+AP����Bk��CG�A�������ZG���{�;=R�ꮗ�l3�O�2E�;���tYg���������O6��������oi	$��a��T��H�Y���������,�p4Ʃ��yĶa�B�X�՜S����O=P{�V���K�<#�������+�8�A�AŞ)	�@��=���V:�i"M\��K3��h�2x2�X(>'+~�w�Y��QZ@-u������/Sd4�܏/��@�P�O\�(��
J�o��=�K�yM��l>�)�+G�^���^�8y���vN8R'�����J��_��((!e��%}����}�I[�B`!=+��?4#���<,��~�N6�D�	��v�>�*�T����Ь�>	��'�9 [�O��:_;�&��㚿#�/z�7s���{cc�j�����h��i��jl��_��RW��{0�G�z~��A�Z�Φ��x�W8xSp��Ԅ�g��2��O@q��J�x��D�*<*�V�U&�{\b���s\^��H-��5�5�X�Bf�8�{O�Z9�'R఩��*(Vӣ͖��r�>|��$W�]1�y����r+4�h%c��+�	[��8�n�46j�ݛX)mP�؇��K��8�(@O�oB�y�\��^�3:�W��@�-9�;�Gh�^�98$�^kRj�%��-4C�9�*%_��{ڇ9tFs�E�	5�r��u��)���n�F4��Os��h�T!��Ȩ���-�]�5�����e�~s҂/�7[q����O���y�,�����CG�$�_�I:������2Q��<�j�.'ނ�c���q�}�e>��%�(M�"�ު�hݬ��((ҩ�˻8��"BݐmV�Ӱ���dz�A�-��߫_�j��~	�Q&�Vi�V�V_�7�M�D��FL�?�q6���%�%�sC�8�㰂����r��l�+Ӫ��4_RR�G���VT���%����6���|�_��[���4&F���H�%Z��Y���qN��8<���mZ�{h(o�`]�UN�Yq��&V�Y~�ڔ�~�VK����7�* l��!�y������eKד�G�>�P��b��,�z�IV�hT�G2� U�� ki�OF�ނጕ�G�K$"ozr1Q^5H7�n�p���n����7� �mK�$���Tlj2�	�|$�
l{#�_ÜCt�FX�0	GD���;�@�p�N�VhF/\����l!���}��R��Xyk�8s)�v�F�3%��-t�d+�D��ApX�Kq�\���k|8��#%e�R�ӦY�CzR/�q��oE��H���FQ8L3�1ZS��K0���-�I�X0o=PA<��3r�X�ȹ-���0�a�5؅����j>W���IAu{��� ��2��Vt��4���.�,�\�6��<�?��%��ʣ	���0�Cr��]S��ʓ��C��H�<��S�����\yL]p�YN�!�b������@�I���;�/�f�Q^��Zޕ��H�}��!#*��x�Cde2�w��KE���S���7���Z� �}�k���±�gTV�̭�<@�=VG`Y+U���wM��%�C��!-��D���v"j�� "M����hDK�m�V�O�tz>�~����s�t��$*X!��ۧ�7�~oE��h14z7��n-������F���e�e^E�bP��2�I�ԓ<�:��n�N���Iݏt=`���nv&�K�7-�K�Qok�H�:ѯk��ĳj�N��s�2+�x�X,�U,=9ɔ��.��d�jX�-}����:k"��FG�&���J�mc��8L��W�.��(M�	���>H�%��w�%�߉�'v+&�Ťu�k�m�~9�=p1z.I�w�qC�mguao%-��������D��H,;i��(ؤ��z���v�u5y[n.���M���Y|8�&j��6��s���|�$�-ƺG�&�6�3.]��n-�͇�����?>��Ē.z��@x���n����ڽ`�[J��n>��/3j>�jK ?���T�yN �яNU&·�ؠ)�Y��W���q�ܓg���QvB��r-w�޲�CR���U����	q��+�=�DN���?���}���I7���6r����I���=��2M���u�A{��Sz�S�y�s ,J#'�b��
j?K�Os.n`�JP`Nz�>7.�5Bs�"��h�J:u�--�"禱=lk�Ѹn�(<��*��FO���ž+�Q�[�|?����\�S����{��+7��NW��8w�ʉz'L�<r��L����J�Y�DÄ��7r�a2!���(>�%�dC���f5)KgY�S�<��(����ޞ�]��i`��O}1c�d����v0���M�d�/�Ch��o��J��E)� ,��B?��F�����E5k��4`��3�,�*=����ر����L�3	t{kk��~y��%V�n�����Hh��h��_˹@�Sǒ��?��/�������kCI�)����c4�t���_�hNï�;m�`޶5�>;�B켾�o�rvh���x2�g���FK��f^�b"�G����צ\vF�Sg��B������2�C2�geː3����q_���w��������%��wo�9��9g�� �}f�n2�A�ޛ���v�#���-I l���R�ӟ؄%�3n	nY���F��̥�����)lq�g�a�i�_􎤓4�k����`?�vbu�Ҍ�X�
(���g��ъ~�� �>�T�G�N�*A{ΐ�]����h�`��#��K5�H�Ź�ɗ�2�������EĹ�X���W�~�]SH�6J� *�U\�y��g�8�����m�O��͖ל>2�{�G~t@-5�]��[�!1�={�w�<g��d�M��=�������b�_4r3��]"�b֎E���y�^vo��0;q�G���Z�7���dp�-[uQ�Oټi����4%K��!�S���� xi=~�
?�w �
H�$=GMΟ�jv�IЉ�?�t���O��U���n;$ɲԃ%}���]�RF��H�����x�9�I� ��pі�� #K8gm�Je�%�_��g(+\x{��窸\��0���/,>V�h��d��4e�� bfn�I�[D���X3�<R�D�P`^���� ��1����[�ҟo�
Ԉ���:�mā���%�M�:2+�:�W�QB��KD��(Lun���H��-��BM2j&3Q�.��1l�^WJ�P�c�&�?D�b/d�-G���kï��Y��5�@��5�5������=z���C �^αR�Ҹ4�g��9�g5�ۡ��E�U왶m~�p;�.�V���yR�Ƣ�T�y��\]�[E��ɇƱ;!Q����h'�$�ס<�qÐjuu���G���`����$�e�X���	^k[%�_C��h��<� ϧ=xݧ�����-C�L�^̨�C�\�<���^/E��;�c�~�_��jvֲ��;&*�]Lx��l$B�8��!�~	����K#��hOo!5���wZx�� @w!n1oy�ZV��<�;@�כ�OW5w�#]fE&e������`Z_���Sa{RU�4b�]������$J�R�<Z�治J��(�Kw^J&a����J�'�.Z�h��Ժ���K�(OrՖ�����i���Į����o���յ�����/5�M.ht�cƊ(�m��r�Yx�`b	��2O��(2�2�/bcQ4{#��k5Pu�)�o��O�E2+�1���4"��?ʨR;\��>o�R�o�	r��s��b-��p��QB��"� �3��Ŗ�C��{� p;��\����h��Vbꀣ��[����ͧ�W	�C����^6�C�G`�!B�y�E!.i�_Zc�*~�ET�׃%�����"&<~�!;�PY�~<3w�t�t�|$�<<E��<J��,K�aSG����� �q�^�qM���_J�9J�fɉ��^�S`p����<)�w�����^�7Q�ʾhQ*J\�EV1�B�Q6����<��D�Y��o2c�}C�Oi��-y{h���%�5ڍ��;\ �{(�12�Y�@�(�C֘�{��^�v��h���R����%� o��X._?>m�V&�'���g��"�n^ߗN6�$�ЇH.y��!J�����P�,����Mnt���EӞ��O^i����B�	��9�31�~�
E�,�B�x��I��q�$g���fkd�*���Ÿx��T�D{J�:�r���bhq��7�86Ƙ�o��cc'�\�
(��M�`�i��I�.�0���A`��w��R�T ��k�f�O4�$p��_ȉu#�`��P:Ifh�A��f�;X&,�a��
'�4�H��i�Eyr��(�s5~Zm��3'I�.-E��H9ǟ^H�v2􍂤���x�OV��ى'@���i��E�`�WH�'W=t����Q�a��Tj<
S�p��M�T��"o%3�i��AZ�d�+!8̳Qk�pr����4-�?O�^\�����	7!r8ddeN0u�ٌ�OZ�@g�x|r<5;�`�����}1Y��	�9��A<��R�_��e@{p��el���T7�h�F��@�f�s��SG��� ���m7Y�����-�l��3Yb<���0�A�ý��I;#�Ev����u^�rLk�~�����JI��쟧���N	5�9��0k�� /9԰(����i��h����i�-�� ��A�G���y7�\z�l��`�.Kr�v�U��<сEz�noyhz;\���B�o��Nۨ��L��X?�����;};�e���*������3��b�4Z.��9]Ä=,V۔��Gqx��-��e�ѰWo�ozi��q��(tS�J07��X�X�d�=I�.`�J��w\��4߷��tT�D?���U(���L�+��@�Ɓ���Ѹ}�1��5����&��Dò}��r`�2���vb�~΍�І�h�C�o�$�5�r�]�GN-=7c�W�ʨ�]k��Y�_�^�ζ�'P'|�����ȣa�s�P�vf��-Ƴ��h�vo-����z��).���؜�H�,��RWq��H�j�V�P�H��/�}M��X������|�iJ�L�<] ��Z��1*�P��c-�-��:�q%��`�ݭ���t�;������-fL�*	�Da+^�%ٹ\��a{�0��8����J���!H_f�
�i���==�g����/��:!Z޸�^����ޞW�e�i���5!��ݜ�,z�f��4-�����n�]���l^���~�~�P���L�kCV/+���wF<2&ל�bq4��s�L�<$aH=�`��}2~�6n�	���,k��S�Hⵎ��N! Q��a@��L�[��V��'6��-�� ˧�X��*��ԢWPy^٧""�j�)Aq���94��:g�R-�D�|�-���Ɏ�7�\{�۳&�~z�i0�����M���sk�bA�s����|`���ΐlWk��C�����U�_�Q/�$K k�C=���I^ͦ���
yl:�R9B�ĉ61o7#��V��v����˓���r��IH'~B%�Y*��yx^�M�౬ҍ�[��U9[#u���0�V��Q@[�c�x�#"ލIT��-�x�+���.(/8jዒ�y��'�Q�!�R2����J�-� �72��e_�ӳ�pЂ�!�\�]`{�8n�k6�?�������Ţ��)�O&�R�\%�p׽��]�+�}�c����Չ��x'���~wd�D2�-�\��KT���n�0j�)�/`�c���I�ԫ�X��u\����m�RUno��lu;zv%zRc��f~t+�b΂\0�?��>�<)�w�8S=LXP����Ζ��5�%�5��(�`����zс�8�Vj5��n#���9l��0������Y���"̈�P�ٮ?i����'?�W5��L2�*��°���;�-ӯ%���I�5�w�t�\�򙿲h`D\�C��"��L��ɦ>��]�5��w�zZ���&r�����Q��I˴Z\p�����i����2���f�|�d����@D\�ֆj��zs�+���'�7ϯ�2V�Z<���._-�����Ⱦ`xE5�Dt�T�ĉH�Rz��`b��҇hv��F?�8(���Wפ�;����r>���M��� �,�/�D���색bDp4���J�ag|�w.�2D���3���S��
�H�~�千]d� ��M�p�N�S��)w�^���'�f��k�o̐��8���&��^��|�k���O�>J5���{�U^��(!*f]` UP�W��u�| .{f�j��xIUL��q�&&/B&5@S����M�9
�u��ݐ<���#�D��|=Ѕ$ �� �`�pzD�J4���f�j͂���n�lc�������/Z���S�|�*D��S�jw�\��Zw�5�W*�37f���P.Z!��*����i�2��;ܓ+��<1���Cf逤�֏͡R"��U�0�Ar��T4'�ͨ�-?du���*�4dA!&�̜:F��vJy��w���{i�Z��K5�Iv(�4Zjѕ�3]{ˢ��Db�;�׍���ƻ�B3&z��P�c�'3�� d(ZQ�=��[�2;^�ӕŪ�J�\��Uw)�za;��"��GSKҀj[���M�0ν�9�A�� D�ON
s�T�/i�Y��d�'�nL�
�PW	n�����,�Ʒ<1)����O9Z��eoE̯�J�ߵ�Ǿ�C^����p�PRZ>}���g20rY�ܢ0�n��Mqi7�k݃�jf×~>͘,}W[��Y'bP���٪���ڗ���s��K��UC#䫘_vo�9Ct�l�|��Xe ����,t
H�j�����5��+))��10�� R̍[�8�#�,w�g���=W��1�E��A�T�%ze@���\��Ux�bZ��K�p��i>�����жL�J*;pc�l��cQS���J��Q�o�=g7�D�틇�\������dX_��યD���1a�yH����Ј�D�`���~�T{H�6`�]3^T^��rj>o��Wo����`,�⡮ KK7�;n�3�説�h}��Ta�dQe���4qY+��=�{.!��N��)F��~ݒ�T�97ͪǥ�ִ��6.�s�./��#�Kcy���2d�gu_B&����;G��d�釗� bƔ]�cO3�Z��L}⪗���2L,�L*g��O�ܭnm$�P\�Lzs��������އ��9M˾��7̿���T����|��)��ij3��ȩi	���S�������u�v;LP��. <����Yؓ[��W�ۙ���:B/�\zl}C�x���	�,VX -� 0��;�euŹ�����5i����0C��լ���.��]Y���m�?��4��N�R'|]R�=K:OMZ��"_�i�]�`�������P�"��o�?��âi1c��yhl~Ԝ�P&mK���\պ�Z�Cͽ���4잤X��I�t�R""�8�g[[L��Y>�T��HuD���_�dx"ȇ��)���2����O(���t�m,�7�HL�J��e1�ȉy�n�o/�:˖�٧2'�L���մ���j��U�PT\�4�|�I4�����'2��y\{F��z�rw}�T���Zգ��(���gz<-q�`�ҿ��<��,��;��9 �?
t.�c�J�d�[�R����+���V�9���R�j}�R+s��ޒj�r��9{���z'�8--��W�b-����������0�s�F&��� �Iw����GAO�鍰n�i	����sA�_5Q������$����E��Ŷ���K�B��	��S.�'��I-$��"���_.���:U����[�F��D�6	������Z���Ƌ}j�C�@�ޠEYx�k��qk���>L bR�+�
U[�36O�B�fxХ��qZ�Hg���ب��4j;3�O��mP�J�D���߳y�P�
���*'�==�8�����)x6�¥&fj����a�<� Zwݣ���ܱ�[����:���޺/%���2��<�#]��$�ƣ �	eءZ���Dar�:��!^���;�`
�������k��C8�te;>?'U��K��M�}�mѫ��X5w>)������k�1-��d��׬�^l���i�W���bU���y�0f(��T㟎Ъ �HM@]m���"���%��!�W��~�K��j����1����rG2$����3�f	r;P;�*[6D�ݮ���D3{_�%xN�!�s��0Yo��a�u�$�ņw@�(�k�=�c��w$�̎���ۓ`[�>�����2z�_�n����їIGb��
�n�����a7��v��>"�N��γ�9�3�5VOKo�6�
G�oX#[��!s��Q�P��#�]ұy�2o����
�4]w%�r�
=�5�0��V�2������2Č2W�u�9]�����V�EΝyO��L��m�H]�ف��g��N���{4΃uj��&J,"�T��$'Q��͹'�:x�6�3ѽ��L+�c��rQ�J����a���`��ut�c�F��T[��a���#4xO��a��Ԗ�f��;����m1��Zb�͌����S��
�+ą����;��ezW3�q���|K�I*u)k5�2����Ĕ������77��0!F���
�ZȌ��v�f�=.9�`��z��&K�tM�~φv��E&����k�᳭�]6����+�@٭	�9�/�5hl��w��������Q��2~i��J�yo��_���� ��yv̒������cuw�ƣQ�+��2���e1'�	��L����y�0p^ ������{����x�,"ΐQ+٘���w�d�#�g��q�l���i��c��x�̚�uQ�m䆂�{��/�����KD������R]�ҜK;�14���������Z�w�g��i&�o��n+��%kC������_�ɲ�,;{#[�egZ`�m�y؁�B�ڴRB�i+���с�.V���"���r�2yC�c?^�8�y*qP�"D@�.��RA���/95P	QWfb���v�z@O��ϚtYgi��p%߀w�6�J�GM��WHrU�o˖��g�.癨���&����`�1�mT�B��a�"�~���7��2�B�W�����㎷�ӕ*{�9��Zd՞�?�w�b]&IKtڸ��y�i��>�#^.b�=Æb"� �O�I� l���<�D���vc�(1���x�b		Y��=_��B{����C��Ζ38�ʙ(-+Z���/�Y���wp�8�?�\���3Ϫ�'�n���Y7��'e�i�>rV"�q�l �RTGk�jz�>���V�3��;�%]��lx�N3�?<�@�>�tj>C�|YOZb��ןEFv�9fF���l�L�t��SR�jО�^�%ktw�0㮩�Fc�0���$�a.luk�2Җ)3����{m��	����?���<-)���ɏ��
]8����O�%9��2�PlIa�$�]ק�썇x����~� ��/���(A��N���Ž�hx������d�:�bk97]�h�?�9 �<i.qCE�sy����Ń�J�lC��ڜ���ɺ�=���7�|D�}0�s��D�\��q�1�@o�/x�� u:��D��:7 |�,�	�k��$��{��6���0�n�N���JA̑ğ���=�,�����?�.5��,$Q�͔�!�:�z����H��H��Fi���~��b	��#L�[,%|�����q��j�f�$�ߣ���uY��#,u�q�m���K(t�hnֻ&�ګ^��[����DT�|�U����/����:r���K��6`"���z���*n|�m�
��¦f�`�f]X�ި�^z��
O=�gB������j3�^qI�O�?j��.��}�5}!K/E�5b�P*�l�Rn*Ś�eY[��&�!�%��J��B��!|�5���fE,�Ͽ�� �1��Ɠ�b�썔�\m�I}.���)��:p��hˆ'��L�&A�̾�)j	���st������&���*q��O���U&�L��m�	?!�1��W�H�S�!�t�9Za�mC�G�x�A(�,]��_GdD�钛�2�_z\�ʉ��%dSXS!+��2����Pt&<��B�|.06%LIR�������K?MA�$��n�Կ�����\#c_I��<�qw�I!`@)cB�Fr�8!kM�
�5�i�^9=N`;
S�ةr��cw�m׸<<�Y��%�P_poG�UŌ���4��W�5���eԫ��%	̉���sl�P!wđ� D�å��6�Z������"��ԟ�Ϙy�!���q
�N�J�Tx�P�v^ﺖt�K%�<F�
�e��TK���'���Lp1B�џ�|�� ��! �޵%U�c����5�E*���I����-�έpڷ#�$buȓd�.��H��4h�y��IU�.=:�(�4D�biTb��~�m���k����^��T*0x��Npo��b��� �F��<��Q��o?�S�������Q�	Q}Ւ��)5@q�ZI�n�eJ��SrD����H74��`
 <���WFm�aTa$���!��'�`��1��8��05�2a8o:�^��w����s������;�`�h�������"�]"N�Drj^|�fͻ`����J�9,V�QG������xG�� j�oc�E�Q�� ]_3��Y�
�Q���(�U����8N�5�����$�[ ��9�1ғƧR*��)p��E\4�h�P�Y&�]���4E�}�+ٍ�F����w!�S(n��C����`R�����Ȍ8��.�/������d�[�mf�Fj��V�ӭ�	RŦRQ7�Y9DN���-��y��P��	A��+n��'r�O�=���� �e�	�"�
u0����ȼ���Va��s����G:Rҩ v�h,af�r�e�F�͍e�NȌ�EU��2'�������h��;u"�F���ɓ�B�	ܔ��:6�"���zh��"4�i�reK~6o9��v$� �S�Sx��u
t]E�\��x��F�����\�'ي��`1~���+�l���"!����M*}W�:�A�!���9I�Y�[��:|rD	=�bK�������І e��L�� �}� ���DK����s;,�LZ�����C�����<��	,�%�k��fn�Z��?�ޗ�M���V��
*B��T
-{�h��z@�W<���׳�!�+Y���9�X<졒���0t���ם&�Z<Gz��W���ڟ-_�i������}/����#8��v�m��W.R�2��g�����)�J�Be�s+�ᰭ����[^����a�Y�L��~�)WwU��`1���ID��s_ �ϲ�Λ�2l
]u�������>��Z��H�]�g=�dZkE���{�t�K0�oܽ��K� �r�⎰�7+�[@X7��;�7���^�{���y]n��}�u6�5*+̗C�ݥաC�[�n�Aa����l5�T�K�����"�p<EC4;[m�+)dv!�ȁ�f�̍�FjR��9J24>�l���w�ֱ^$����h���5
�"Xx�h���\F��jgӾ�'� H�����L	�'c����G�\��A���K�D��1{JxlU��9�P_�Od����dΤ��]�k�w
��š	�������f����K:
hq�E��Q��|([9���0	�O�A�s�F�if� ��3Ӭ|E'��g�Sͷψ$@B\�\��G��ӡ�ר�#��R8�/�5�e��q�2+�.�u�P$@u-�Xb��U�4�{?�I�,	� ��=x�_��q�s2�J���M6F��AT�Ml)G�m���]���Q�⿩]}��,\0��Csr���i��q�9�cw
6�b|��(��E���*�?��;^F�A�y��;�h��ݬ��:/ivA���4
P^n>����y��~���~-�o����&ר���(C8k��v�<��դ֨K��Z`�#K�\R���Ά��m���lP��$��R!xI�e�a7E����)J���I����o�6�IC��0��f6�H� �WW��4�"!j�軲���� �`<�i�+��
9���uzg�>����/�+��|,J��X�w���xkd�N�k��:�Z�Yz���{��,�;��Ʃ'�z���#�*e�%)�RM3��SI��Ւ�8��q��_�{d"��a������QFk�o٨��w���!�b�MsG��m��gͻIi�!c@G�"��c� L�X½�䜨�@��O�v��c�)�7���d&B%o������usA��0�(�(����>_�����f�"���(����L��Gd��J���ʓ� ~�/W�����b�>4EnGY1�!PUV	.9L�~=��9C��N�]���d	�S��
���V�`S������!#�RW�/�A�Ah�7�u@�z�T��`'�/���9ݍ�(/+�W)�`3�͐^�NƜ&jnZM�w[|h6����z��i�i�_3���9����%e��8~�X���F��Ik5������p�̄`���a��o6�(.z4�A
P$�i'�?�,�����������Ն{ے�6�_1��vXԨl��O�G=�r������}T�6k�Wڀף�F�	�j��o���h5mcVMd��Bf@$�>���ڬ���൥�WD::�����C�s�����o�< ,��X����$˟-����4�r�׫�n�`����h03�;9i$��]��*�<!ٺ����#������ʌy]NK�!���e?���]k;��\B����s^��x�"��ߵs��{�놟�Yщ�\\��71D%��%�N�]s���Q��(+��蠌b�眡����Lg�y�FPJњ
S��\��9]�`�Q>&L(�j7�t���?t:rK����h���s�#B��r�'���ll�#�Ӱ�/bт��4�}\މ;syb������3U�2��e�P�E��s��67� #|&(cS ����ξ� XJ}�`��p_��M N����H���Ud^*DwƑ��+(޲<�L�S'��x5_-;Z��L��T���c{��կ�����]�6�.�+0�|��S��\+puiN��+ф%^����"��$&"��Ӎ���dsγڥ���L���_{��f.+�|!�����Wf�	b4��_F�0t�l�W���/�n�����k�P��L.[�������ǥ�
��\��s�C�fj��L	��M�2��GGg�m�7�[���J+`����(�	��d�L��v�SM ���Z�_ْ��BI,:��H�V��ommɩ��u@3�+L�Au�Qŏ�ԥ�ui)�yZ,��Sf��
�<a�M�c;.�����<g#=12�]Cq����*�z�N/��D����m#�T�<+���,�	l�U� v,�iMd�ݬV �%��8��Y�bY�h`a@%����'X[`�WI�G߸�u�n�
#���F-��ޤ�Ő�mW��!��Fù�����q���w�-�=�}	iyz�*v����ݙ��k	�5S80O�/}�j��������>�g�S��^^8�Z}.�NR����V@
������f8s���^#ޏ9��\B���>���{i��t:Hx`�v8�{�e'��և�I�,�P4�����]Q�w� ���;�^��MR8�GVt���2�]�`�R���B��o��7Y=��e�_S��F^{턡C�L�~�3h8
��G6���#$���[`4"�~%#ʫ��p|�U��N�GӪ�o��5��}��wd)X���B�UB�_����×"�
�Y7.��yta��d��6[�f%����%�x�X�Q#p,�O�A������,��,D��2vm����Ur4�G�
u{Bת����%)����w����CZ�;K� �����=ި��3<�t1����-8�&Pw��<2d��� {!
�v�×��#Z-��U�X̦/��_��=���EO���W�20��pb�6?��)X�lE�I.�����&6�1�C)����{D�U���1X���1�c`Р*�4nf���芿^��gB �D��%��� ��r��'�Я���B#��!�"Y��>�k>���̍g��c0N�2dM���䝔��#���T��Z�w:��7��&ނ�mut�c�ңd�ξ�e+,��h��5�J4��O�$���Prq�_߼.K���5&Ch��&����Tt;�:H��0Tc�N��Ba��d?e�_�8W�_9���i4p^�j.)����^�aBc�Kr�s��%�^x7|��f�����
y����6Z�������8Y{r�{!E�ND���v�"�D�{��6cϘ�S(��)V��h�80�5U�µ�J9�[|M�U�e��m1�.�t7�]�f�Gu+�"$��_#]���^�K��f[�_e��0+.l�|��9�ɾb���u��6���D�IN��;��Gk�<f���5`���O�F(	�0V������B,��u��5+�Y���E��ZovDSgm���t��#v:�ϐ�v(:4�	�]a�E -�mg-V3M[�0����7�F��_I�8E����05�io4��<eU�������H���6�,oKjr��G�.m�B�B��w�&�Uu1�U�6.����������bŰ �1�z
v+6�}�L��=1ќ���/(8	G��=���7Z�*Y�7No$�m���&~F��͈���`��m�V�U �`��s�Y�:6-n������e��H�{�vGS�0��֪����vQ6'�H�6{)����X�fr�r��%�y��L?*;��o��>2>m��ِ��������]z�| ����co*���K��s�:���A�0r�4����
s����pU���<�o���B���\���7d���N6R�k�Fn*�9����k�@�vk��Jqe@ų{��d�"k#o�ٗ��J��-���OX{Z�B��c2V���˅�G�#��m��N��eT6ɧx���6�[��q�n���<�(q#����������Gf~�U�u�`��}�G��T������r��$���N ��̐�u+�A��pH)<��j�jݚ�Q���&�K��N�Tx�[͋�Pc�H���چ�'�xUȫ�:�c�u`Z�ج� �,�v�c,�!�ĸ���?�i�;�{�ہ�Q�aN��O���j�J��Bp���E�`(N-g�0w*�yVy��I�BjX�N�E9.��w�X�TW�ߘ�;���|g:������/�Mmp�"	rMYX�╫����G�;$��A8M(�������=y$m4��-YɸñV&�"	����O%eLS'"ő<��>�&&���"$��|�?�f��J��� Ч鐃C߂;ЮA������F�8��c�	c;�M⦣�A����!���,,B�l�a���#`]�v2G�-�4�Y]��<�%��ٴ�8��
@:�=�m/T��ܠ*J��vʱ�.�uU���_U݄���<V��n|~���^�]D��x���A�P5����o z��=���9j�>�O�H��m��<>��h���dv`�/)%dJf����vν3$t�*�c�r�����k/��J���k|f�V�*�HW�;�5�%�I��-��v/�2�ZK�vW@�L��U�(���,���17V��gS�X�D-}���yS) �  g����],$��Kl����iQ�9^�)!�%;��_��1���2�"u��kL}=���	vص��>s=���E�Nb��.��A�k�~ҝ��m��_�%��U�%!h�5�d�_��%��r���s��P�<@R�t%�6�6V�EYv����=�����&��8ki�F�i��㻮������$�~z걁��y��b,���OT�������H�2JH���g�羺*�_��/A]@�~�3Az���K��(�_.?JECL�{۸!�{6��/p�?�]Q w�@���M��`�{�V�]T�v�	��bc�����V�32��_É�.E��0кT��˘�k=�C���il[pk� �LK0:��=���z>пU�d�������Sc-eQ��;����Kv
�6ea	:��$B)íe5A{C7J= ��ha\��"��1I5����]��钍n��)��!>SOX�q��w(~��p�F{f�wh�\J��r��fs{��aE�۫E�@J�y��G� 5����~�%��M:a�-y�I�jWT�C�	����cc��n+��^�5'q��i�3U�}�� ��h���Q0���m��`��b9�/��C N�	;Z�r;&����/�-�5�5���ұ~��Y5ih�z�0��>m�,l�O/}M\w:�By�kfP�Y��H�n����u\pr��]rtD�����$�Ԉs�:zT�ʯ*�zU4�֧����n��s���
s����Z�Ix���D�֚c�צ�U�g�t��=��\�;{�����1`����s�/~	��Q�q�݉_�3oV+I�����G�ԃo���������}�}c�nq�. \X��0�薚��S"d)�ć�+u�P/�NW�9�E.��6���B�<QE����Ǣ��:�
\�"����~�"�x\��ܖl� ���y����j���1`j�=�(�&m�j�>n:ФV%%|ǰ����cE�� ST�|CrjQ����]���zL����Q�`9������d<]���;�S=c�%��Kg�U;F8K����?�^3%��2��̗�*�5�@�T3k
NL�C/k�s�d�x��7��a��gXu��;E���xù��%��E�t���B=�:3��v$C7���]��I2�`��Q��A.�ڬ����3.,�8����-�mSw�ŹL�q@-aB7���k��� ���{��[7�f�$�*D�rV�����)�:9���u�}��.X�F��mn�R��-1���Z�&iE\` 'B����\M �5	�';��6i;���H�9oXBN��_���3�q�a�7�-��I�/(�[�;�y:>]-(n�vE�Y�_��3���@UT��>���jsQ��F�#5D-�>�D��*8���b��' C����Č�-㤓����4ف�$��@��T�Q�e�8�E�#7����n��<S|�aGy�&|:�xG���u��Hh����#-H��1�0~��qe6/�wz�r������WR����3|E?�����������L��'��ga��l��gAj��)Ӄ�NlY�c���ꔴ��DU�Ĺoa+�0�wA���MV��������<[O}���$��T_��(��X��cﳱ��H��Z�����c����K@����[��ܶ(�د����d9r1g~�C�����e<)�r���F�ڪH�N�=�p6:�I�l݉@��&PMF�v�J������{ɽ�������Lw��P21�\��vYMM�0:��4k���s���Mf��a���J��"sdT�K.������u��K���oNݰ���kB)`dc���
�)��1�	?�nȥ]��I��,��\��� y�N��%5���1K/��q�e�}+��N|��z�R��67e"4����%~t�W� B+rY�a$x�{���~���/ 7<�1�[ę��'�W���|�&X8��]�*�ǝ�g�n'+Ln�E�ˡ�#�g�g�x_�;�n�����e��o�W�R��sp�R��W6S)�G�ڼ�m��/�eo�_z��7�J�����=�iݽ?��\�U�������}.��/��#����
���꧗"7n�*R�	A���M�FG+=t�>�Fd�b�8��T٣�MO3���~�c�8M�z��Uh'7fr��s��	�-�E-3��|}'�o�So�:���������g�[Wa�AI�2ËsL&4��
�u�}�{~K�`����>�~�7C�xW5��wm�c�ꉣZ�1K��N{2��\m�R��(�t����W����g���/��z��ԐMA��װVd�e�ۑ<��z��D��,�Qj�k`�C�^���FY*��M�P��N.�?ſ->r�]T�+)�xDT�Y�y|
%�c�͋a+@'NX��Jt_���Nkϫ'��2�%��/b�/��E��;V��{��b5VrbD���0jQ?P��M5�m���N��d�3��+�݃8�9}�.�F0�Q�pQ����]����yG�3���9�?��d�0j
p�v�O��[Q���<��6�[���gO��������𡝸۝Z�6�s���p�d�����M7ctT�YP�̡�S�#��G�U�?�8���z��Щ��ӓ�/?t:�+��μV�3Ꙛf�J�L8Vp���uo�wę��	�fw���o0S[FT�B���m��r9i��#u�酴�g4X���*1���A����͕o��~�E���ΚZ��I�q+BI'���1�cQȃ~� ]S�\o�7-��-GQ����M�X������C���ߝ�n�r,:�U�^p0'3	r.�M&�~O��'��R*�}�S��A��B�0��M�����E)uWQ�d!]6�C�n6,H��F�O�����^���
��[��Y �R�gk0;��*�e��a�a�WA�4�h}՜�y��?~�E�:Qf��e������k�̩�C�|
��D�ד�`��Y\YGSe=y�ώH`gDQB�l����@�P`<�P���~�G�&G�C�L�X���-�G;�J��5	ׂ^A`������x�;Y� �q3�p��`k�ٜuu�NY�[X`Os��5��.kt�,�M�VvK�-��Np`�Io�ov�1[ϝ�I�s$DD��BS�s�(��'�s���ټs�R$�jO&\�@���v�R���a��>F��� R���j����|JH-u���yA\'|���/*��k|UW{t�[D�R�G��^�7�61���?e�8�U�ܯ�M��J�#A�-t�x/nz���Z�=S�<�\~����:5���_��|R=��q���������3h�����.t�.JR�қK�w��[�WA�?�~�qx�bh��"B��;ٻ�b��X�zp��ݶU����t�K.��)<@W�k�.�۔�/�����D��@�+�A�d���я�34`����!��_���zX$�f���Mӵ�������6���v�����:��d�������T���9&��Ι��	
�g��;%��M���Ǝ���}�/E���@�m��Ɣi5�To�/���e�[�9yk78|�Cy�Z��UT�H�\5/܏L�6-�L6��5�Ϳt��&��5
��E�ĄG8�eC�j�x��_Th�L��A��S�?��JU����q���=f�o��>��,/�=�� ?��_���=���@ĪNT�K`ɣ
�e�/q�g��u:zDn2�A����ژ�jK^8��w�H�/��-|�B�7��[�n��}DD�YlĬ�+�{�DX;��*z�49���-�D�R��1��V��Qy���/m2�)D�qD�cv6}{��rjHw��&�� ���+���_˫Qߠ)z��>L�C�L�(�V��l˝�����N��܄��<'�EX�a�}�p�����@��-Ȼt�ց|�w����#��gV�wn/��:R�2��������hv�4��`Mo��р�H`��W��|���RtO��V�W&il����~?���]N�#�g���C]��<���[.�0]�W3��د����q�\[-.(�=I�}�9 ���ŀb�W�1OߑrlQL�4~�c�Wn��21~�`=�|ũ"�yz��rU���qZSVo���Kڼ$�%R�U6���l5�F�S�8���O�"O`^�y��1(�;�K��O!�Ū�;Gis@z-�h�2h�w��W^ �����J���F[F0�g��>�,�x��_4%�3�˄�Ir�c_���B�5[RO0�)h?�W��ڪg�m��Ύ���JOfl|TW�&J��I,!�_ʣ��2�״ԟTQ�}��Se6��1},y���I?�\H���͇C��U���l#���Ό�Ɍ9".%il\��<��-F�Aߖf�1 ����A��4zA���POK�Y-$�G)����j���_d��� �����V��_�&�1�A����^a����5U�闩�87����򏦪��	�?a@XХB,#���ZL�r��L�3ll�p�6P�q���n�=fK�ܚH���lX�� 5�A���7��i3)��u�oG����,gT�ح!�#s��5-'����W.-�f����3������e�����R��4�5׼z��Y�il�3���'h�E��]��	��Y@����=~�0�X���*�E뒱*w�]y�����{� ���|��D_O@�T;��L�����z�O{������Mjq�ʰ�R�e���B�Q�d <��Q���A���2Z�-��o5o&(ly�tx��ȾI	�D^�����Bu� �/D��g$���$`���6�/����VHPww�=u��cA:>�T��X��P���dF7�ڄ~���-o�����:��l+���!��/}�jX}f����u�R��}���dޝ'���i����W�;�s��,�]��ү��y�[��}q�a��GW,�'�~�e�s5�(�-�|}���-�O�;۱�>�;�0��W�_'VQ�b���"�T鹋~��T�kF4����^m�G|��"�\�%F�=��xW��\�]��v�,ܬx0e�Z�W�A����	���E�
��_��OZ��h9�V\^I�Kc�Yr/�[�*;�`(t�.�8kȾ�{�e61�ٛN��ِQ~�`D�#���[�����Ż�gk�\�.�e\P�)���)r�K��41���b�_�T[.�\�z�R��L�H��P3X-r#2�>�*z]69S�W���� �M� ��u^�%�����m� �g�)\X�!���/p���(@�4���3�T��i���	�M����㒻�V��ܢ`%*<%��i�o������¹)z�o�ϱ(���:��e�S#��%���EX�*�tp����?�<�Og�I�m��^�c�kiV�:��Ȝ�u���ei���0�����5�;�jv_�Ďm�?��$��I���ΰ2�(����=yg�g�>��d��BF��[�{.�6���lm4���F�K��uh���������
%Ad��ʆ�G����h�Xm_ri�G�GI�CYAk���� 3�r]��RV�]��7M���wlR��BI8�	8�K;+U�ӑ�go�ma��No����<��w��^�(�����^4*M���Z����vf�E�
VJ6��Vp���s��\"zn�����BW����iE�V:��^5
��Z��	u��H��\��W�4�no���� �D���o2ĦF� �G.��F[��0�)���|�q:>���,k��;x�_�DiK�2�QW^O.����5�@@�Y0�=�H��|P�S�WD,����G�ݛji��b7��]������K���6{k����Pq{q!#�Zk�?w���b�7k-�o)��C;=���S!Q�q���*Ó�N����c=��֍ֺ�E?�h{Đ�f�/�sMj��R��a��g���� ?�¢#f
Y�%[��̔�n��`���W[�ȯ�)�\t4���54O׆�����h�}���ʚt�x���ig=�T��

6b]��h�N-�Lj�[a����?�{)r�jʡCg���j��mp˵�e�#�Ua�R�O d�fo�ڥ��h;&�8v�,�hv؉��jӔ��ZK����T��j�$e���ڶN�!�ޑn�� 7�������UW �M]�d�Ҽ���]51p�#}�z�"��������x�I�C�f�Ss��&�|R��!J���%9i��(�U�^݄;��+���)_%���6���|�m ��x�@�E6٠�*7�N��:��{��� �P��YJ�?�*��J?���YZJ�����|���p�	J,�h�MտW#_M	�X�>�"8{ÓV���>lY�����l��� ����G�ߩU\m+2-ǋ�$g@�f�^�f�ImӅ�B����r�ſ�]��`(��	_�����%$��^W�X+��7�H�?�oPb]}>E�ᠫ�A�EQ�7��s�g7ك�X����D)�}�ޟ�	��� z�j�Ph֔���x��=�S����<]vLs��L7��(u�z���&^;����v'9���W�a�K�:]ΐ�.�
B�
�v�����1�;n�
���8�jh�����(�0�~H.��P&|�1y�Ao��9��A�U��H�g��b�9�}�7l��+W� wӺʨ|K����x_u�O�b�� &q�>@�T����;�b��_!��C3`���h*9���?Z8s�4r{!���&�ƪ���7�O!�M����yl���ů����M�)�V�>��:F�`���Ǉ�}Qٻo��gog�?PV]C����1>���&�q<��"m�ƥe�r����ǒF@��]7㕊`E$�I��E[1��k�з&�!�ܴ�N���Ju��t@�ƌ�C�r���`\a� �C�[�S�i8������R^���;�� ���,�:�ӕ�#���v=�ÿ�5.����l���{{�g���A&������_&�������e.�h��f�5�9�&�a��=Y�߼V� HE�L��ژ����#�$���
�z(�o��hr�l)Y�XZ\ZD�9g��x/�S(iu�����/����+��\S������%~[�*V�lc�C�(9�Kʒ�� ܪ$�Ry]&/���(-����<qu�5��_7�?�sW�H���;h-nCyO�(%����{P���Md��eA��F�MWR9���]��J��g�r�f���U}v�~
g��:�M�YY7"P�<��6\'�M���,�p�I�ۭtl�ȑ�dJ�s��*Z�C�9�C�ǿh�ѳx]VO[��9��5V.'�
3 ��!����-B�8�u��{Ɨ���`��S�1p���!fyP0�"��$Q2�$�2q<��K}�aH��ߩ}�I��u��YO9�.����w��DZ�R��庞�.����\9-e�-�����!Y3��a0�<��=>����J��HL����&"&�ϐ��Q^��	~�Lu��<�L�M�� &jo%�Q�$ٕ�[l*��;��+�_��z;�t�?�z	�'�c�0^�p�|H	��6�����Ed���!���$6wcZ��[��5����_�Ӵ�'c��
�c��`{Wt��棱X
u��Ugsc��������.�%�_�0�u9�W<�1g���7Q0�/�c�/u�u��Ɲ��f������3�� %}�>�	�6��n�����ǟ`�8٠���"Ve�k�夬v�����^I�A��YAӷ��3�����ˬ}�W#G!E+l�U)���O�O�D�,���B!��zD�q+t�hw�|h�JʽR�iU˚�R�O-s�q`鄠�M��ıVd��x̑��%�]ߙ��w����BA����C5l:1� �&���h�r���	AC��F�����	
��: ���S�+V���_�p$���h���:����W�@�ǈW��.�����P���S������5%E�h��:b^�|M**��b��J��/,hl{j<�S�ݛ��b��/�0��Z�w۶��h���C0�V6r4��f_�d <��6�7�,��P�}�u#m$2-i@� :JZ���VF�/G�m{�6W-�-8u%g/�l��ZSk7.�X���YVa-���Szo��9T-
kC�_��Nv��RNf�R8K��$~��6��'G�rKȍ��ރ�ު>G�꒣K걪)�������V��Ӊ?�(�t{�`x�զ�	0ޜ��p>~BS�'u@�a���-�ܔ�:p�1�F����V�#:�����~��Q��X�����sa��TJgd��V5����	���[�����������7a�:߆r�i	�YX���/�pT��7�!%oGݑ�p���K�m�;'k�B�~�z���o&W�S}RT�����_��B���zͶF3I�~��(��z�F'�S���$��@��z���w}I��&���c�l�"����+j�Y������b��c���W����Ij���S)	�l�M�wF��R2/E�Qx�0U��˾��r�`]�ֿ��Ѥ�B�����W���D~Іr9�o���//�»~��~(D�����e��M���:��+*?��)�濊��Cp;�6r�
;2�8M�^7 Y�E��y"c_���s�r���U@�.��1/秶^`���y�<}���p�IJ§��j�Oi�me�Xp�����KE�3w�K�!�-�vջ"@�B����/���F?�□�T���1��RLy^ˊ<�`e)���0���� �`�N���
�����TrB�q������ G�ڒ�������U��dR�*彖e�4�XU�1��=��4w��P��	��2#<y��Mn���O��&ߊiȃ�F��*^Uմ)C��'����M�lFtр�zj��.�վM�vv�d1A�q���.�����s��No��,�iw�����o�(+tQ�(�p[�G%��	�"�L)�����J.q���s;��L��zX�kcr�ܼ3@0�}�8%���!�9P4����b`u4B�(��q�	�A�N��wlφ�P]|��e��c�Sy�)Z�V*O]j��/Q��Lp��SF.�����E"<��1%԰S�@���_�]�];{ѽ꽖�%�ZolD�v�\���i��O{�Q�E`����R��ɻlL�r�?W�NF�$��x�����kվ�W�@�wg�W�d�38��юF�e�[K߁���~5�����
I>����)k�s�m��Ȓ.O�)6�SݞtšX��1(��L-��ϖiH=�f��_J��4������f�{SE�Qp�Ѩ;'y1�d�h��W���Mj,uԑ�h���6���ҽ%�!���5.����~����OY�XP�v-g��E�EQx���r�wMߢ�f���S&��۟p��f�xE��3u*A��I0�����N�B��}���Zᮼ��eGrUb�8f�j�p9w�c���{T+~�U��[���ǒ1V��OB]$�`�WT5�h���:=�̃Ҧ���D㫱�ѾZ���&/�v��J���J>ͯH[��c���B���+Kx���{[o�MJ��¿�2u�.p�#ۻ��"9��*�i}�DF�=�'Ea�ތ㇕�{�Н/�9�gpH}d?�(�������
��}>���]6PM6�O�x�hzJI��|&��S�L���ч�4�7�D��S�Xz9�Yu���#g�lV[��5o��I#@DѮ��qsw%E�z-��x�����s��&���T�J*�܆�#[J⥃���%����,����h/���jxw�Bn5��gu����k5��A�����,�m�M1�r��B^��"��19e�_��۝&�eu�Fw#�l0�"���BJ��Τs��l5U������J�Z3u�'n�\_�*�әƈ��ӹ�^�-��V����f-���U׭F�� ��F�ms��A�QG����ҫ�Z�}� �d��|�(v�(�����|9�J�R@��^�y� �#��S�v�O��~&ի� mA2��� �YҚ.&�>����to�����Qm)�+��l��wl{�%�^<��3�-��t�7dY�a�J-z�e�Q��iӳ�����`���Ԯ�s�(��kǿA�;/ŶUj��X�(�����X3���R�Sغ���u��KESϯ�%'���#b���0¦!�>g�3s�M�6���tŧ[��'QXaH=NVj)�
}���A��a7z���N���m��aH%u��# ��l��z�4�z�Sr(}���3��2�g�H}Bs�w�L�W��nθ:|t�:	p	��5]�˟���nW�V��L]E�E�u��(?vAW�J�ǿ���[���P(ͅIVޟ����^({��}f�(g�rg��5��Y�+��;Yd7��s�bu'_zAa�d��7n�.�n������^쟟P�q�m	s�:�@|�,�K��ST���YJ➓I(��u�H��g��7�}�j�c�T	���F�(U�<��F^|`�~��))�"�����Y������!`�\�o�cwvnhx2��-r47{��S�/m���=]j�]���d�%M%)�f�q�O���	I�9�|䆢Md���	�G�M��q3K׋�����e�**�,i-з������f5L�B����ZqxϦۈ�|�'_<u��Z���tR}��}��4�f�ѧ:�Q����8IIJP���f�s����ԳE�N��۷o������ۧ��V;��P�� .��gUd�x`�+���g��\�Vy�x��jN��<o.�~�{`�5��v�'��)d�^Nn>�������8�ݺ��z��٠��~<�)�x�"x���~w��M�5�,tV'«��w)�Uq��-��qp������ �E�t�H��ڼ2�BV=Cѣ"%��L�k}��~���?��:Y~��Y�d!\R�@WƴB;"�㊵�(ʙ��GU�� �Ƌ�B-�7�("�^�q�ɹ/���O�Э��4��r[@�-�pl��RY�Y�X�l�Y���9�Tϥ��Fu�ڶ�ɫ�韺s��݇�+7Q6�*�4�Rh�D���'�nΫ@�.6�x3D`N���4ڪDo�v�5�_��f}��r��ڡ�F�͢���x<?&��T��i�����w��n	bE��pߊ�(�Љ�0��a���)�9a�c�h^��Ч*EH�P;-p_�?�!G2q�K*��4g��&*���I����JT6�?�	�ure��ό2�^�s� ���$����u�x�m�1.1��M%��{�@�k�ɘ���vV��=��?̉��6:�-�"[����Q����C�5ܖ�7�S�"M�(�j��F"��V鞣�5Z���s�
c�*h�Q勿~a� ��{��$�(>.q��ӢC>p������5�����|\�U� ��/���w�J��`X$ 4W�be��L�H��O��9ݜ��k3��^{���L�_j���s����C�(�T��Qӷ0z(��~��U.��nZ\�y ��E�SN������\���x��9B�~��_��f� �V�KQ�js�B���`���2	#��M���
�c�Ë�C�"�1j�5�g��a��|��_Ȃ����h�S݌��/��9�n�V���!D1X1�j7������s���3��>�X��C)� ���=��>u�4�F�{��1e���0�.ɐx��n(�ڠ� |h�c��c�/�J�(=��͵��h>-[���e�L(�Q)�Γ�Sx�G��%�,
2l���tNF̡R�y��W�ֳX4N��}�I���F��p�c��1:	@���RW�*)J���^N�e�Eֻ����^��D��=(��Zf���ѕ96J�"P�|�B�� ���qz�I���[���^�_�B���,����%7B�a˶��*nL���0���#�1�J�o�O�C�yֹ��f.M�q�G3}���R0���4�n�� �[�n/oA<H*�S�1��8Jv㼡h��a\{��n��H���$�l �}l��&� �ۏ?���`��H&�D8��ŭ���}y��{��:��%֫�Z_
����X�6򕁔���*f12���r���uk\x����������Y:�L�x'�R!�~�
A�{Cu	�[eh��qlD�����G!�\��h��.W��C>v`�}���Z�����%���+��1��G�Tb�|RӃr$������B��ۊ癲�l�V��D� �y4R���ٜ+Y?�Y{�5]EX���=�|!�"���_m���N9-��ςTe}�z��'��߿�X�f��%�b�2Ж��1�.�ML��J�\�i3u�u�A�m(+8-<�AA�c6$��֧�����k�$i2�E�|	]%2圛�`=�}/�֕�;U�ϨLm��۲8����:hrJ��.my.���-^ƹ�pi�P�e3�ěOf(�؈r�oa[�_�˟}\-�#O�w��L%��:�D��m)�4�X�gl=@���MAK�0�i��a�������&��u�e���*sZ����O��iaY%^���֝&kg_��N4���*�7i[�;q�y�|�%8��O��S�c�x���C��c�|a\y
 oCJS�SM�����\-"�t�q�6��$�W���!�ˈ���ae��)-	-���c��Pkj��_�WɈ%,[������(:���4�%�2n���p'��,�`�yR�
S��͂U��\��Y�=��L$��Q�UMA9���%0�Ƒ�2�?�3<�IRi }�B	�V�ɴ6s�;;�I�n�,>����,���L�������"����3.�7�F9�䚒!k+	N�!��A��<��:�E�~Cnm?g??�����ٽ�=7�{�l����!0�m�K�
�)��T��S�� �r�B+Qc؀�49�3�"˪��8�am8L��_:�A ��LrH^�h��(`Hy�Z������6�@_s�����:��Ȱp2@�N���i*�\� hXiN.�{����|�v�?�XH���P풴�iǈ�4��+Τ��d6�0|���GH�87~ͨ�o��b�TiΦ�Į��y�m���S��=�8�K
ݶ�|�~\ń�t���(NS��h���;!�V�гdV���q�ڥ��-����������F�� �U��Z�vM�x���#L��w�|&<�����ԏ�,&�5����&}���)�p4~����ܵ/5�\/Mė���"N����U�$���c���7��k����c��j��ؠh�*��Q؀���l��9������ձl�l/R����U[��>��-���=kh7�/j�:X�Y|%6gá���;�5ˮ�;o��?��i�t�{S���D߻t@c�l���c��������Rx��<83M�]��g�v�C�y�//�=��>�4�ss��6�������o&�����ˬ��mgƊ����|
&M%�N��e,�]�*�c7.�ONً��u��@W�M�z�z�ca�����Cr �X�[-�T�
�������<l�M2~���^��*0�/l��D�F�2��$-���JG~��~�.f��Mit�U*�C�P�؍��m��� p PT+m"/]���g�P��\Ѣ8D,���ޟ�p�аY�sx�(dWC��p���YO�fH]2���rNv6�[^������%z.N�_`��Ƈ�..�����O!�;��ç���������1o=H�hL�߉Ag���y$���J[-�(Oƫ4U�1����̙�o(K�G���"�,k9�[IU�|�-�!�� 5[�ϓ6��vd:�C��Uvi�(�&�P���?�5{*��b�r����GW +(������ra&�P�Y�H��?I[]�>zJ�l���D�@O�p5�����	���/��iNh����Mb���HS>�*��
�W�����^!_)�O�˗�l૖���Lr�{��|�{1L�|?�8���dXY�v�p�	�qH�[��F�{T��sJ��~u�x�ċ�p�<�{Dɏ�ȅ�l���'��ԚN�=˵�@r����4��R1�,�K:u�����q��qB��(����y���;��TXhv6����7�.��XV�d;* �P�ыm�|����o�m��U_��#:�5�`�O������W���-�چ$�M�kp�(����>��8��N3�z ��i����a�K�#��$x����I<I�k �?���.'�s��%�`�B�*��n������[G�u6�����E���2j]���-ͷ�����d] �۹��z鏅��C��-��J��?�]H T檲
צҥX��M��r���M��{w�\�����D�9���S��U�<����=�8����6yQD�����TG0���ڃZ��1���3Q�c�n:��!Q�v�#��b���QI��W�_Oy���-���0�nJ�բ��zj�%Q��@���_�`�2���A��&B�& �������ښ!P����@��^���߉����G�����F��E��I����&��n��IӔb�b�]�a4$��z����I,�Fgs�2�R-��a��.�⤨�އM:
�o�Q��5�.���������D2R�L0��zY�g ���Zf�޴�@@�0��5��k��TT5ϻ}����8W����
�"MꞦ q&×Z��]�3x����[K%д�w�m���U2�?�Nn��_�M���p�e�r\ԕ�Wi�#�q�g���w�������3$8ru
�u�8�d�_�z�/K�+Q�M���)|��݇5�f�;�7�b$�VE
��!8��JvsD9�Pb@���B��u$9PΘ_���a�AC(����c"/�����G|�<nS�rG)cԲ.T�/bgk�
ү�N��!1W��U�w@�l��]g��P�7P�"G )|�ᩈ4�J͠���GF�?{b$��N�`�(c2���*�e8�vٻ��zL|#M� �]��$a��'�X7���3����,h�Q>�e��Φ��qy��8�[j�ɺ�$���ߟ������l�9����kW�PP�*sd��K��VB��b��>��NADiW.S�+���J���&s�}_�E�~����+%!s��3�{
6"�;��_s#N�K�� C�(�&����O�� e�=Hp^�(9�[w�N��8K^�셒�_�n�>���z������_��a2Cc�z���̏��H
3G�\*]�O���j��*ݬK��>hKyŭV�gQ�C (�:Z��A 7���{yi�]�]�d��@T���y�o�;��W8@�.��� F�S�婉B���u[���,f��ZCL�'h-�_���cw�K[؏Z�/�`�-o�ƈ�ma�I����e�<nO���Bw�Rl���+Q���)��Gy�>�2L� ꊪ/�!��1QV�+��c�ybL�����c"(�J���z�\����v�2&�{��}R�l0J4��y����TƙQ�����%	��.��^��.5�J�"����&	�bI� �V�x��%(���K�)׷G1�]�ֲ凰6Q*/h�U������E뽵���YoSO(���K��}^���8*�Bz'�'2�i�\�T2���Y�q{�/�}��O�ei��z���FI�~P%f������h߿�x�ƺC7jSÇr��W�\�P��^w�m��v�Qv��A%��F{-&�J��~�@�}����Q�`.�J������";�~�x�<�N�I�x��Їw.��˨o��"bfT3���]b�|/�G!������s_1��7��FYp��{(�RH���M���b(A1� d�1��Q���N�u�!�н{*	�#"��Z=�9�b1(�D�Hc�O�-Ih�yM"����mGs�|�ܵ��iy~���'�l.��	k���Ⱦ�N0�t�x97�<kdG�g���sH��>l��=�h��o�n��]��$۾(�]��Ԩ6,�f��
���x"�o�p�(��0捦�q�qh_�N,�(UTi�趀q�>䡯#O���Ύ�<����5�����25o�wD_'��j���5[o��T���@܊�Lw�)�F��}�G�W~#�3>Q��C�1�]i$g4��y�+�3^�|{ͿfV�aH�t��n���(�+����4��מ�D�]5� 1��3�8X8ɚ�qSlw�-�7<���3��1��dѐ}#��o7�5ȂT*o���2h���������XU^�@�'���d	�Hu2(t�f'�����͒*�At;Ki��L^"'4�[�$ĭ,�( '#+T&�bR����vSٹ7��u�< m| v+q��3'�[+�M�̒�4�`�-�V�Q.�#�����a�\B��p}BLB��R,/?�E0��J��F^s�{��n+.�b6���h�����/��q(="��H|�$�+�y���"5�%@mz���|E� �4@�7丗u"�MQ�����c��� ���� ޾LB�,���R�k �� q�aV'��"���v��m������P�&�'0.��&#]w�F��ϋUE����&T��)$]36�]'���"@��(�]�A���f�d���ɦL2�\�U�?Tg�q�
7��?1��7�)[�Ʋh0)��;4����v�s��x��)4�T�b:t;���rt�������.�{��`&�����vO��L"\��܈W�k�t�,e�Og�ʐ��Q/֗�؞ZŤ�a<�jaT�_|5�ѷ~F�0��޵��f��\>oh7��(�tl3����K�;n	�K���g���/A�t��z��V"����6��
}��h�K7!���OA��cv����\� \�-�ozY�uoQ/��{�OaGl@b�z6���Z��#�CƢ�)scJ�����������o.j�#t���W7��ہ���������Bk\�&���m�JC2�Dj��"��}t_%��k0�q�q�X́�y?��>h L�%��AUp��qd�)���:06�Q3t^������;�:V7<���h��&��gT�=�H� ̂-=SOS0U&9(?I�r��t�p����0��눊�`��.�F?1��$���/���%���`��n�@lVs�_&Dd�/�j�R��Z���Z�)Q�ּ��Ңb�bU��dVZ*��ՓGI�!
�zʃ!Q
�
Y���2��t��<5\x*'��5m vC�d�8���]���k/�Ą�����?]K�����9�o|9�]��9�C���&��V_����\�`NһH�?�*�Z��]Lf�����D߅��������;��n���f���*B��خ:���%�1v�yM���Q����q�D�I0-��j�1�J.)7�����ѕ�jȞ圁��3v9��YS���hƑ_,Ļ��G����nͮ�svX2���C��_�<&ō7�M#j� �&�����s5�|X�՗N۝M�n�
;ZC+�L�@���D��핤Y(˪����}�O�)y��}��X^2 Q�%����A;q������������� �r�pJ�*�i��� رB)�`}z_&���7_Otӑ�)Rnl��#�dK���<c�� A؋hB2`ሩ�ξ���<����:��UzՄ��38G�G|ԫ!�a�Ʃ�z�G�n����6Gh��j4D���ئa�af�̗⠂8�8�G�+�X^A�5�M"]��>�1�۫�:��*�`���S�1���
g�R�E�.E��^�f����t�5��㉅�@<�{C�ء%�c'8C�r+C�-����L�(�4ֻ��vt�IĻxi�&Cl幄/��#٨�w#�e�(��>&���(�����ɔb��׻�Km�s3� ,9*#A�7�$�g�{�ás��(|��j�$�K����W��[��_�+r���>��J�fq���sƷ��X+�s6��G�Z�"��"�&�����ݹ7<�z������.?|
���L��[����j�8��Q18�܀z�]����axE" �m����ÙzT���C�R%}����V^��/�L��ݭ��@�Ď�݊+?I������y�窺��G�k��+���P� 9�ʨ�y�v�Ɨ��+B$��7S&�Ĝ�3L[nfg�LT+�c�C���e2�>)Y%������_Z
H��Y
2:ց����N�_� �vJ�BC�DUM�M̢3k%d��́�4וfDGÉ|0�_�6h��N���xU*��)Y�(OO������3��&�X��Q��邿�O��P�Kb 3������9�mjĠ����;d��{���ۺG1�A��.���,l�9����`+����W}&�y���#xrK�`��DR�hkPf�__�dn�㕅�-[�X�9ԓn�X��	�rY'��\�	�8eZ+�z/�GR�%����K��6TR��~��T�!jJ�d���xB[#+������m�]#Gɀ�9�}Iq|-<�	_�Ô~�xl���Z�k|V�f�uX�������t�h'+�Ƿg �wU����՚OF�(�YV�h�� \��B�\��mc|���z�@Mx
�-w ���U��l�E�9������Zu�1$�8��s-��u5��m�CR�����h��� �TvHI<��a"�ԡ.#�w��7d�0]4'A��kn��Ֆ�N�<me��Ј����q��aC"0hH.�z�d�˳�1�i��%��ĭIvf�!@�}c'�m��,P����(�g��wF��#�AKp��<���}�U���^����it��ݹ�SJ�2 ��mV��I�3f����t��l�y���>B�O�+�h�+�E�8�5ȳ�(�M�]�EǍ��e >���쭀2 ��v��co���quKdk�^�s����=��g�9�9N��F@-�&;Ez���z�]��@F��Yy�e�,�.]�X�1����v�z�w5��-���o�/NΜ��{�k��=t�	3���0�D����2/�0�@|*K�4�{|���h��4�k�;�U+���,7��a�D�*-��2i��zI	�:��?����f��=K�9Fd� �R8������'��4��%1_���@��xb�R��<^���8�Y$cY�㌽�fA\>ID�Z˙�	�5��!T�CۇVV�� ?߰�4!�l�1�� j���7�јc����aoƙ��t�8��d/�yL�Z{0�p�
�?�&H�|�إ-��N⯪���쨅��+lSę������ �*z݌��=���H|]��[�ī!�ꮁug�����2H�s���ڋۘh��Xپ��c6)�R�zbh���bu�:Ɓ����ء��������ބNO҅(�z}�ց6���慏�{dE��HG�8�]���'��*����{Kug',�pb�t��3�^�"�xz���X\:��ɒ�k��VL�|̕�,���ɜ�g�r�iݔA:�oj��r�n�^����Q>���0(l��������ͼ�ޞ��'�6&lϱ�o��ИZ}����Fp����eN�2�����ox�#aZ���_@�^q6��3�MZ�~�,4SBX?��W��:VcrX�������Q� 9�KJD�wr�tp�'��N�F@�]���?��v�+�Ǵp��G�H���Y)��C��B��v���\5�'��WF7�T��t��Y�'��v=d��ui�A�/���7�8j�-���FIk��rJ��W��ѻv/��L .b>�� \/1�"(��m���f�j_�@_�؂�5�KS��4u��1t�Ľ��!x�g"leɁ$h�#�x;�9�6�-���V?�M��{�sb�����E�ٴ�E��,���WV������Ũ���3�ZH:a�_��f���d���ӣ���/0� \���9b
)r�R�����+1+�35�[�/Bm*;�%��s�8��eyB�ye��Y0i�ܧM�����1b.u9⇃3yAS�����@�&�J&���C
�GՖ�?9��[{�ޑ�0���4��'`�)�f�Ho��Ő��/׉P�6+F�k� �cl��~������u����z�B���Đ9>����4���2ċA�I��9���o�k�9��+�s�S"�M��<��|��HWy�~ڷ؛%�
�fucx{���*bÃ�kq�M��^�oK�{c�y���?��l�b�O�0MJOÀv�Ɖ���/3�h^FW�Y��Ն�� �O�6��m\�\�6���8x�3��\�?�'�{�u8��챨J&?����':�����wzS�f3�X_3���	�\�_y��/���L��\;�zBx��G�h��:��M^��$_)0��S�>f�"/���gb�u�r S1�֚v��1�[?( ��%So(#)j-��઎u�-G�3�����d]-�Mڰ�*�P���������O�������7�������寧���,���Y]����]�Z��6�4��;�]\�;�Ђ�zR1��։��̆Z<`ͭj��Ù��%׀��j��<e�0�MU���9o�'�
{��x'	�/඾�xp$J�<|4n��)okt�r``�1Y�ݵK�����+`F��Ǹv�rǂNQ�ӎ̲�4�I7S���Ov�������ec#�M����.�I���s"N46C5�ih���e�F�����,���۠�W�)_l	L9aF�ny��~�%��0��d6�����MK!q
	�2<"v���s�aOL~�9��v��y~��fŠq]�%���cv���I���\�C�������-)�f�X��>Z�	%���������s��2�I5A����[�~E/��Ǽ0�:rX#X'�	l�<}t`kF����G�=�lД ��`{�a��1��]H�t�߷���w5���T�xba2k��W�̺	��������tKO�]�Q����:����{����7��[�j��,���#𞔍OZն�u�!���Nq ���$��J�}
Ny�����?�l��9"���߁6��?��&���>���[/��o��k]�y��H�t�mmE?��g��F��9��s/����M
ݙ�L�aY#�����Ŀ��l�P�O�����)f^:�?��b�O��00rٮy�C�׌����Ш1�ə�)"��h�sִG�)S��^)��h���XV^he���^����`���E��=Ka��dØ1������ߌ�K@?�VLS��r�.s�{w��~pC�	oN�Rk�NIzk�����E КU��]���6���X	2l��z��T�.O��Ǘ�1���z��B�����I�w��������ꍺ�o4Mb���tJ�tYol�D
A
�fV�����Jm�
������9����� �!�b�����R!,�_ŌHlvAx+��# rÜ��k�wz�Eƺd/�������)3/�GjU9jK�N.v�g�<̉Ȉ����42o�B׏h�<M�Q���x�	�Ol�(��=��H&&��R�@��5K��(À��A�I���p�~\�*�Ͽ�R�S�����̵N�|���	>�i�4�B�a`�������qX���
cwкz�?V������Re�p/"����[�I�.X�Mf�Ge8в/��R�!�aL��X\`�	r� �A2�F"�=����
Ԛg=x}�%��lJV��/�M�T�ݧN�G
*X@�� �͉	����5�U�<&]D�-k�w[0k��ps��aP;�24Q������.Iܤ$Ք-�[҉�H�@�y�s��L"n�7U�%����h2����;4�2�w�c8��x��չ��ۅ���9p,�/�#T�&<3>$Xb�����,���Ƨ�z����R�C�c��,	��-~�<U�U��ؘ��{%���;�s�x� j+�O��NuNSxA3$�6	�B�
w{��������-ϟ��E2����y������K���:����������=v�Hn�bO�ĀA|�k"����Ɯ
{`�~���P�����/��*]�_��!g����aA�î �R���aN�E�H�'mA%�j������J ]t����,
"�;H:{l̩���A�-���
�KqTuOb/)8|i��)���	�+�0#x�ITFe0]���e�1����_�C|��o�ح;���S�D��&���!_Q����	��V�P��ڽ���L3[���ZX��MӇZ��I�k3T�������	� ��9����Lj!Ľ����rbi)���t
�D�al��8���kP`�.��H����~P����R�僫
�W
�!��p卵F�8/+#%�$��Z��Qw}���(��Ii�E3��q+x	��yA�u�n�6�P+-�O�3�[�ǛT �)Ä�Pv������P�"�6�؈�GK�Xn� �M�Lu�+�zG����8������芋�
%���]}��_-��XI�͖�%b���8���Sk4�s��v��5Ω 0��=	����U�F���8<���^��.]c�����Ӷ�A���Mz��z5���?���9^1O��H*^q	�Qh�!�g�I�1�,���c)�ECJ��Ƃ~�y��NDr"�p|��ŭQ��ѭǛ�c��2�j㮷,�����,Z�m���Ո����>S�y�[	{@�ˡ��O�Z����#�����S�w����N;�/���D�i��Yыi���&%��:U�6O?�􋅊h|�|��o���i�HC ���X.Oˑ���?39E�й�'B���X;ְQ\'�y�:�������O�p��A1k�o�{���Y㡉�ΈN��X�*��\�d�;_�4ȯ7v]�k���P ����a
:�M׈�-3�	P�k�f��x�GT�s� �؟~7ۖ�E
��:II��M���I���]��(�`F���ޖ���K7�8JՉs��<��*�K�0,�t�M�N��iO��ְr`�"��Pn-~�
"���u�Z�q�����hV�2�P숬��k�Ln��U�/�Q޾��Z&��G��'~�<R7�(�X�H=*��[i"�y*��*Ϳt����K��b�:���ǎ}�{8(��J��e(7�X�$�h7x�@|n�F2=[����� ���B�x>M���T^�û�	CD;a]�EČ)�0Ɛo/��Z�]�{��%�iX|8JH5��lDY�$Z*9�,�zk⁴��ĵl��I"7�eTq�( ��A�='Ɇȉ�)�V7`{�e���;A�lҢD�������:�4�U<[Գ����y����¹�M��~�i^oD\�!��0O��@����2LŃjî_�e��v4��C���˳Jy٣���I]6�	���)�1����w��#���X�m�ε.�*�^�QZ��*�}��I�G�H
���̫������o���V�z5�+Ĕho���H��:>��{pU�(#'N���=y�i�@��N�3M��șM��k��n���Fu�?~Ҽ��PZf���j��J�{Կ><�*�_�V{r�m�']���s�B�@B;5y�֕��4��\w�|��68��,�w�dy�۰<��}fI󅨄�x�[�ײ+�����;c�7��x�kr��]�]����:Km���&.OSSɘ������):})����
/�؍�!�*�NVvT�,�t��*EԌ��1�3��<�=���WvX	�A��*$�ج`>>����%6`�� �&U��FeDM.PƏ��ly:4򑘚�P�Z��K�TKsO��(ń9���M��d�vk��i9���L8X�#?�@�2tP�)]Ȕ[U�$)$;8��S� �I�!���J������¡}Bw�[������,�N�<��6Q�l,HD�ɮ�HȵR��y�^��9eC���s=u'y��N�ؼ_�(+�Hi��%IA�.M���׺��PjP~���N�6l昮E �K
����^(Uh%E�Z����G=�%L��s���N}�W �G�}���&5/l���<�w�b���Θ$���a�:KU���g���"P%�%R�׼��Q�tPi�'g��X��E�O��X�Χ�x"�09��p��b�IMa�j'ި���57
;��A�Y|�B`Mko�������S �y���)oxR�A�����^���o�:JV��^ ��a�����K�Q�d��=M��
��T�I+b}DڒwC\�-�3䅋q�*��ά �ȔĹ�Nf3|�R��=�#6�ȴտ+~�9�P�l�;�QP��Ǟ�\Z��5�M�	�6�V5o�p���Q�_���>�.�la�x�91	�WХ�+3b!���q(� =��"�6{ڏ^�������ff�� `=BN��$��.�.�DP����`��!z��K�"�~���PѬ�eW��D�^��	����G�E Z{R�԰)q$���ڸ�q~w�@�w ��xϮtX�G���-�qe�`QxX���aQ�� 8�Lbs�������cs)�'a���#S�jh6)Ai�P5��g��v��\p���~���̇+E�9_���|_�~Imk��؋��o=ߞ{7NA��}�=<�u�Y���b&́e𩤹�qPkҘ�Ҽ�x���,�n�����i�_��h_�*�]�n��������o�Q��SԢJs��lkVЋ/@�4t�cMA���v�����'��b��W�8.C���W䈑.�ġ{a1����=����O�����$���Mo&	���l 'gl�(�*E��B'�;�k��Dܮݙd�[F'G?�*�����������kQ.Zǃ<�K�w�k������DV�?��0��ZTt'͇Ɉ0h4B�IyJ'�c�Zn�+��'zP�{��ߴu��цV|Y��f֭�[0M��IQu�/�)�ALTΜ3%=rյ0�h�B����wJ�:�~b�ai��^�z"�=��0��m���rV�&�Uw��2�{�"�N:���/v���}��>f�{Nv�U�t嫠7�����,�6�WN1��0<�>�8��`��	���Bl|�,���l�����Ĭϧ,��Wj����wf�B8R���wW ���5�H�}I����v_��6�D�U#~��8ڕ��7� "J�����]��Bi��>�8_A��G�.�m��Z�
��k>&���=f²���n��p8]���$4�8H��]�\#�f��S�܎�حO�{�3����8�d!�듵5� ���T�<i릤}�JKY�+>P���\��C���7C�~}��F��>ظ�o�Xu�Tz��V�qPw0�Vu��j͈��?qؾȴR �X��aD(�R؟�:�d��'�u��7^A�J�ܘ�$�q{R�xaƝQ�z,��xDU�es���
Y�Z��U��(�[�X�cj��PAw��c`�	@��(��S/��~Y�C�Ȋ��=%aX�f��%2��v��*x+��/�{}���M{E�e	���C9�}�̎��1$���vv��&�K�]LYɫG���0���R	�����A�Ѿ��V��*�d\|g!q%��Mm�*'�������uU�C�~d�kS?���0���7�©�;�,x+"Ѥ�Ua���ӛ�sP��2,��=	�^!���}�"��
���
n�����WI�ON?�699䛇Cܨ����h	n���+U·Bt����,|RC�V1�˅>�bw*��y�������7k�� <Ǣ4���'��5���P�Dƶ#���<�г1�dX'H�%����/w��%	0y[P�G{�hr��r���,w	�)ߋ5Yξ�q�\1�7�D�D���-�+�T!�֒F>H˼��A�Ur�K><�V� ��l�J"�c��uaL�EUD�@J�v ���}�a03���������r�OW!���!|�,X�ᦫz궑���qD�.Es��)R
ӫf���3�t�ᕑDօ���f
� !=n��ON�ˮ�pt5�H�!o	�D3��>���x�4U�*/�>�"��~�#I���p�ݏs�3�˲U���Uv9Uy�.FڱF��o�tIS����O�����!�7���!ɛ�5G����m`( i���F�Q��%cȿ�ii��[(ww��P��@u�>,�q��a�ִ�6�F h�X�ca�;#�-���U��R�wQl� �!��?�j|�����f����_Z����~�'��7o�C:I��2,���o��z5��*� �G!R���=~�����ѝ��-|w�8�-0�I��K}�=��A�t��\r�P�^�6@T��#�eA|�k�E#Ka�ܵ�#�� �F�U����xL'��DG^�j�1]6��]��E��2�@�b��0>L0u�j-a�lD<��oIA�.�S$(.RT<�E�*�vd��c~�먖b6�^�D}a��Ƞg(��Nf�����C $�`�C�����*j��
�%Ǭ�2�m(��l;����8���ά�BT��&��?6�F�H�!�{E a��s�h��_�A��o��jt�X�U�7x������,k"�����t�7>T�ҏ�&�a�$�}{ֳ�6^7�v|�P9��1�z	k� ��;�ρ��#w+�,]� n^�]�ǍJ{Σ�\��MN/T��LA�=�t����#�y���Pne�[s�r���1P�L^�?WYk���ݗ#� ����]�eh��K�?>��e��%�׍��3�e�ސi6�� ��PJzm
*����y�<$~���������wV�9�)l�/��"	����6��j<'z]�|N[��\	{異d�X+�l���k�[�/ �(1G���?q�/�i R+nA�O�4�\Xp�{�(wDu�?�P�?蝥_���&�7������K�����%�T�A��J�����rIm��o)I��v��Z\>�Å�z��*���<)F]9Qbz���@P�3q�N�H��T027�ҵaݎ��&�1>���ƮG��v{<2�-��O��5�pUf��<�E�G�b��ϒw?��g����A�%�7����(d�?�|55��r�5�|�#��s.AT��n8��4m�BA~��*�s����9gw(�}�&�V
�0��c�I`*�d'�Ұ�1�z��������AV��?�\m#g��Ôp��s�n��WJ�G��4 �4�F"u��*��T��q=&, 	�����I{hx�	F8 �r��h�����U���!��2	&�H�kb(�ʓ�ti���&�zÙN���JK:����h!�m-�$*[�W�Ds����6ڲ��(T���G�1��^�G;�{�Kئ.������&.��I�n�5A�y�6���J{�/ź7LM��i�#�Ct⣇5�NO��7
�z/�$.8�DH�-f���;�/����\�WXlA�,�s�r/6�[���næ�ȑY9��`C��c��YO�1{�:̇�%f* �)qr��_����=}�]o��N���^f����>L�>�ܳ��Kv�u�����B�w���d����;zK�b����o[�q�u=>4��sTt�G
���#l�웷��܃+H�IB9�&�0��A�a�����$`���)����{�݉峵�Wx��m��llo��(�w��������a{���.��Ws�l9".���l��Vw�G�rwAwv%��e�\c�u�������&NT j�p�Z����컯�h���.�cE�f`�q��/���>�4���U	Y�	9�%K?U��9B�,bt�s^�XW�ڮ���#���FX�+R���� Q�4�����pt�(!g͹�~�}W��7n��uKԫ˻���M�Vކ�t$��S��~>�1�R�znr�@/���̢Z �f��U���g7C�&I�S�E}��챗�`Շ��*gi?T�-�vS���$��K:�i�ytQ%�1�SA�;G)]�cM`H�/�9l�;�=m���j���ɂ�'�:R~�����ˬ��k8�!D]G=K�|���M�j�������˕�bd�G^f\*�IUl	��g���]'�t��UI��X"0Z^��2�C�t���!/�,��O)�K��.�QQ���p�WFׯ��v��l*�\�)Τ��e��1��j�������H�X�RP5�L["|�PG���)�V�dA��^��IT�I�P��Țs=�A�60 ���*d	�q�,[��ݑ1@����(z6 �&�q��g>j�P ��3¶�8��������C�zcMQ��6�e=�1Lyȯ�'�J~� ������D����{�����5=Ng!!G��d�6��fn&�M�k�u�zB�,��"V�Kz�,n)�U���h�Ѳ�bĺY�םmͯ��gG��7NM���\z���۾nJk0jI�X@G|tUpʠ���J����3�Zb�W��l�z[1��[��Ĕ�  ���m5{�N c�7�A�`)��W�0L����:N��������  ~�'�P���ɲ�J�������Y��ҙ����(�?|���g\�I���_$j$�}>�O���RDIۯ!�!4a��ﴻ����f�΃3���u0ޯ��'؃#fc���KH�lӠ�M��y�үM���{�z��L�>3�u�)��1*�J��{$��xJ�^}�S].�Y�Ds  �䙸�?(�-������pW���|��B�_�4���ܪ!��7�6����I��T�L���;��ƯO�V�!3�o��iLV�-����p�+<r�c��Z��N��D��mE`��~m���'9�f�J�_����߉	M&�� ��?MM����QH��ui���S׹��C+.��M��ϸ6����[���oV�R�y(��G:��	�[/�S��p������(�1��;ˈ����E�;%�tǞ�1͝d���Ð\����@a��x��W0�lBY&�B�spl5l�����Ɖ-g2��?���j��Y�X'�Eڥ�K6[y4�ۜ��:zQ�E��=!cx2��p��-���M�^�T���A�Ɠ7�,z�b�*�JC�� �#�~Z��;2d�1r�.$�X�!y.��z@/�,��P,�	���袧
, �d�,&]��j�&���sl�lg�v��C\�"޾��(4�q�yZY����m.��v�d 1���<c�0f�+����SWs#_�q[x#�l���ȁi:ɭE��Ybmz��4��^�W��nc� W�9~���E�ۛ`ؼ]�u}v�f�:�� ��Ow!3�^+Z�I�>��g�(���5x���v|�77�Z3!�H��`�傶�3MD�W{��>ys��͟Z,B��/�+`T���?�l�
�\G�Tz�]�;)	��*��샏�-�\�
�������%�����x�g��4�d��6��q�!�ꂍA�!�td}��6�/=��V����Ш��}�#�%��D�tz��!��H�� �T��m�)�������K�4�Y*̄�.2`V4.�jMM��?Z�3�6�g�zE_���J\��血��a�Im�I�Z8de<W ��B���Y-G�Ef�C8?c	&1!�vy�`���}(j�ݥ2�.Ӣ�9�X��Uk�v�TL�Jc���w�B���L?(�FmH�,,�d���D$�*�Q?�3��kY�v�'L��F9����wo�M8.
H	��ú����@*X���
T���s�G;���������]�� �u1����`�ꠝXP�Y�l��_Ŵ'  =�5�o~+x#�P�V�� �x �����'����\ʓ����Z�0���+s?>;\�＜��D[�c�_��^nXG6����\�H�g��]�Y�ul)D�1Z�����_j���,��ή�<UU�۶� �}��=���#5��^���P�789��檛��
�ׯ���/�.\=���â�����
�A��i�R2��pVQcG.�X��\�}�������"�s�NPyh`'�,o2�4��ky� ��SG5��@1�go]v�N`��;��O���8sH��q�߂|E���R6�ug`�b��}�T��:��ឣ�䛊�{��47�����0�a+.��B��Y�_:F?��K|t�<ר�BV	,ʅ��I���k.���L)˨�"�3�#����V���vV����������{�G��nҘ26�Ƀ�{��j%q�G{�N�����ɭ��$�|Bsl�*��+�3x�`�C>�W�Ss�˒����h[�^Q�Q��8�p� ��d<kһ ����:�Yy�I��3)�&��C��4��\ᗲ�#�E��&~�c_+P=���ӧ瞊�=<Q�{l��O,��|�mUU���@�7�ܴ0V�T�ѿ?��:��D�`X��h���%���"�O�����͚�2H~��(�"�\��|~�#�j�G���������S�5���m"xحo�Ԃ�K�b��y/e^�,	�F�J�L���}8kM�7��v'�6UI7E�Q5`�XB޺�h7L�*�m�E�QGF���m�F�&�&d<�>K������͡�c���qfԖk�2��=F�����u�p���k蚇��|�F�E��B#��p���}L��z�%��j�W�| ��n��+�!D�>I��.V^n��RK��7&
�ms���޶��w?��Z6��j�=6c��2�b���^%���N�FF�����4u=� @f{�����9��]ƀ�D,�[Jl;��e�/nA�)!�l�1�J�+��#��m�A�-�řL �lRY"���	��B�]j��Q���$kF(�"���p�4���X`���Za�
`���1l�b��~x���LYɟ7#�*�VR����O�k�`����/�Ŀ�J;F ��qh������P*㶕�f�=�2��:�>��:�▇��B�,t�ď��`�ꁫ����I+��A�y!¦LR,���r�q�'O<���Q�m�B_^{z{�Cox`���3Az�Z��Sy���+F��,�!Ȑ^��S���V���j�͞Cm��5!�*�;��wt�[خ����
�K��D�Z�'h�2jU�Ɍ\.>��A�F<6k5g�'���",��������!�GH�NɈ��x� G���2;�o�v�����|�&bU�<��^��W��T�Jǳ�{�Gt��w��4(F��%��(���&'���'Х����9��EP��K�d�M��z9��P��yp�K�bA	�mu��������&W��v�gF2z8-v+�+�����%˺���3���u���F����X1�!W��w���4WL~��D�"i�s�d��F/E/�x+!/��Q6�D�8��L���۔ӕ��	��E]����MB��z����X�Y������1:y���	��:M���5v,� �pܞGLe�B@�9J��YǡMt>`�Z�}RX�ZRV&\��'����@�ס�+��乾���l`g��%H���ܻl�򖡱H;���kI�Z�/3o�����%K]��I�
�/r�hH5 ԙ�Cel���*[l��~Y��B�B�n���V )�A�*�{��
 �⁵p�sk Q�^Wg*�̇����lk`��ı8�pC��y�W�Z�
�hd�8>lɄ�r�*w�0���vc���BP�0�;ǩ���lUC����[��JA��L�n�:��x@*؀�2��=Q�^��rR��1Kl
���!���������N�J)>���i_>:�Q�`�(���Y�岠VܦI`Yݪ���O_DG!^�@��7lm�b��Hl �{�
�p�f�Y�is���Ϊ��]�nnn?�'Z��?7 83�e�SϺ�}�Y>1���j����ڳk�:DA�O�*t	����L_x� `�/��!�c<�-��9����6N/"p�ٻ�^M��h���.�FOa}
[#�v�X�fM�z�
�we��Mڀ��E=��$
)S�B�$�'�c���<�߽���Х��e�A�etfG�_��m9L<q�"�^ʝy�R��4,�%�}򟹽v��#nD�W�-��V͢5lĩXj���6�\�OW켙��E��g�|#8�z/�\E7�R�x�~���n��E����Y�cgJF�}��'8��E����5Ԙ�\!zek�>bg�&Nv���T����|f|�0}��!.�G��5~�_x���آ�Qn�ϱ�-ÆM��)l*KaV��.���E� ̾3
���~�j����Yw����j#q���Q�����*)pU�|�p�����X�m�6]��(!E�K��JXr'�x�^�������M�OVjIY���:���3"-��@A"e��3�r���O1j��+ �8l�d��]de�ҌL�HO�@?�wTš�*��k�0���̨����1�@�.uW����>s�JH�cn�l�ӘR���b��m�B�p;���R����Ϩl�c�P�U�A��uaa���Z$M>[4��������*�R����z�m}*V�����{�V�YGbj�c�	:l��*�sArl�.�?�2���*�l����N�Ig��ެ6���q�t�F�9�ya������:(�[����[�/�y[�4�9�>��=դ��|���~�E���:ԃ`*�,�2tF��V#�c��9��^��׫��J�Xe�m$d����zd�		��'�hJ��$`�u$��RgI�2F=;��Q��P�cZ�i�U���
�F�&����lm�C 'м�A������)�4�w�.Z��H.�q��S�H� L���
�����h�]5��d���aַLwӐ�y�A�t7 �T�٠6x�B�C���c���Z�z<9��l�&�A�e�8C�	A�zk��Ȇ>���D��Gx��w
��s�O�hK�h(�O�J��ѝ�"[dI��*l�x%��O����c��|{�b���%:�;I�g�ԍ!����ʊ�A��m��%�ե�b�j���&���8�V�"OH�2�a������h��7�
7��9�q�}�qe^ �YJ��k��+=�a�^�z��7 wl8@���Qm��	P� �%�k�BD�����x��~u��<��5�	Sb��]1�t&�qpM)�أ����\0[�٨��6�jUX����~fAE~��n�Q�Y���gߴr�y}ur��;�Ȯv���l��e��D��"�]r����DBE&�� �N�����ò��-/c3���+����ߖT=�ڑ��)�{��!�Ʃ�0��t?K���7��s�]�I�D<]�$-�>u�l�V���i��6��ϧ�y��R0���ЧPX�ߙn�ۦ�09x�Y0�V�X瓛����x��W�C��n�_lC7*��QW�i���qc����V�h��3�H��P�ƞokyll�[:�?F��L!?p�s>�S�>d��T���=�]Sj��v���o�zLx��~9>��I���lMX=�ۍ�^L�1�>�]�O���:
�{%8?���9̡��q.Mr��^��-��BԳ��l'{�/>o��+�k�QFV�5m嫩_\�(B�]�c|��c��<��	��gD��/���.��H��Jq5�O���t#u_ *�r���
\DA�����Db����Seh�������S�7��/�|6�Ԕ�A*��Q�SБ[C��A�����*i	,ѱܖ�aV�U}֩L�?�?�'��xm��T�O�t���l ]�+�Y�
p����J���A�Q��핦��u������@��֙A������j�����^��qàS�
�	L�B��]qJQ'0ڿ�H�)�=I��H����
���x�G��=���-�	w�A��_uA)�	%o�Σ��bJ�i�u�R�&�ָ�'_�̧~�x��� Z?1QW'$��cvnO�@O�p�|
|�jIRvf�\���m�%�NղP��, G���>��P&Q3d�Si��7V��J��V��c�őuj�Y�?��*&>S�5�pw&�2ҷ��p@8/@�s���
�� ��S��20D�y��+��4r�i�M�s��9?f���*(>4��;���l
��rￕ���{� ��Z*ؼZ��$4�	�Ix�LJt4"��pSτ'��6�T�ƽ*;m<�v�O�׎����~L)ayN��Xh�~	e'$�#,�*�0#�;��Τڏ�����sw͇iUٵ�e-�ѻ�I�F��GQ�Q�f艿&%p<iى�����+�U:��
�R���S`\q�@�]� ?B}s�*-��1M��>H
�m,Q������C�n3����
���"�+cRz�Q�'�I{�nT�^rIV"p��F��,���?�K3Z���!�tiC�H�)I�q2�H��/����1�Y�"�ۿ�=U.d���=uhK�g�g��xA*�%��,Vԝ�;�僧r�[@k�1y ��� ���7.�zO�f��
�&�S Eh�e+��N�:�p�L�>�3�hXT�W��Zb��Z���~�����_�%�z���W&U����c��tB���\"B�
���v�fba�3�.@���??��i�.U��u���j�Ϧ��!���p�l�>�P��@��/�s�^��u�r��]��aqю���z�r�%K,v8����� ��]
��d�PW+�y���,e޳�<�;���D7/iN��{O��@�f�ߴ;G4��&HS���d袳�/�r�(y�ܰ�`$]��^��"x9n֍q0�Z�f=����o��C�(������	�Ik>�{���.�R$r�S�p�<`q��#��6�
�%y� �:c��P����鼄���~ ������X[�b�x[L���l�n����ă�a�)�-g����H���(��I�a��R����F���aohl��;�d�4YF�f���
��r��/)M%�h�����tʜ���xmֺd�x�T���")�������5�``iT��N��� ���l�@�<��)�����0��K�,E�_��v�=��⒯��s|�@1�W��RO��؄�MŁ}�ųUIgp�������Y�14��7Ě���ۭp���`P+�������yG��WC���(UZm[�Mr|T�i<*�}��1��/̔ݽ9Lf�Z�	T�R����N��Cjn��I��P7�\�J�~�ZE���1ׂtN��u�.�ſ�|q7���h������W�`澲	����jTW���H�E��:(����JU5�{��i���D͓��%9��K6�y�:����r�HT�dy��C��p�#LުM���e:�b��-$f�^��x�t�}�i�:��%��C
^W�@Iܐ⍕��-��b-iCE�ky����"}��1	�i4Ƞ�:}'
�E7���O~7҃z��06��ik.�\:ʪ
Ņ� ����
�[��d&lq70����Z9=��3���'� _~5�x�j#[~��q����[�u@�_9��#}B#�L���7����wc\-���%!(^�徾���
�_�����9D�����\��g�?
�|b���"zB' ��T}z�Z�S��y���C�y6b8 9J�#��.c�a��H����*]" ��Dqy�	z�����/���X>�Cm�+��������P���
��9=��[�As�<���?�oa�`��ۦ�/U�oY�^������c�����w��D�7���)�t,��z�'�iV�Z��������~�u������"�P��Q��z����)=#O�SJq�2̰ќޖ0�-�\�2��W��6�hn)�d�����Z߳�`�-�=S��W�;�x5��KD���$������zqJ,���ܯ �Q���F�<��Ƀ�d͵vR�z������ͽ�1.��p����xj��M�2i�� �� D�N]�d�³w�@G��^J᠟D{Д�䜭��wk��nGR8kH��ҡ���*	�s�BK�v_�d�ּ�,E��E���3���6� ��,s�^\���o�� ���vO�U�>��R��i�a��.�t~@���<9|�T��A��6V�p��|FNV�C Q��^,�]?V_��|\P����W����{%�htE�k�o���K|�u��:+���G7_�x����2,tS�vQ�؎e:Ұ����@�|��#{�Z|��a)�-��7�P�Q���
�ďZ�j�;����O�R��_r�`���&B}];�X��oޫ�o�]7mR]���G� ���Y�(���`~�nґ�m�Q]����Hi}�>�d(y�Yg^�J�ԕ��ɮb�P«�gM������=Ǆ8Xǻ�1���)[���� �{s��������C��q�&А�h]6��,�����Q�jgFnޗ?xᓆ[�[��%W��T�Vh��c���)̘є�}�"�@�P�2b�BU�>ˀ��	;|� ����dL#`��xЧ��=��9�}����'�YF��7�l���B)1h�&��Z<�����m'ͤ�8n���vHb�V0�HN�=IԢ�ԍul�"Z����K¥G@���p i�i�}M�#^�<f*n�4�j����|�.�<ET%��`Z@��腘� ��P�$1����ܕ�u¤~�+(�Y�X���Zb΋�������}��Y�6JBd�q)Yu��m���f����yb�s�$G#�T�B�5�;�Wa��%B�W������e���t��;/ԕv�|#�[��L��%�ՆH�����ڣ:�I(.'}P����˙���*�*�o���^�s!����ä�y��(�!%�;T�vW��	R�L�bw���B~?�d�<�\��������������V�D-b��A�����Y��*�"������m;�WE/�xC3��|����$Q��yX�~`�=}��h��W�z�����EZ���O>d��z�2wI�:S���o�e������8 ����ٵ.��E�~��܊�� �Y<)����h����ܩ5�-��rp�8�6A�����E'� ^�|-%e�D�)i#s��ȀaPn����{H\GS��J��Do	E��Ӗ|�5*�;u8vC�/c�>9Jb2�{���Mc��Qy�_|t��������wmϢrz�S#rw	!���6Vf[����ʉ��k��:�B�mZv�!�Y��]�S^�� �yɸ��R,k����,0 S��[~�KI��c.hU��V)�f
r��N��
�-�V�uɰ0��˽�@]?�;(�_������8b���&����51��t%2Ĉ6��]�\1�`��J�?�����q��DJ/j���d�x���%�����(�o"0@i/�WGէC���RG�3vے3q�w�c�� ��Zg^�U<�߹�M�L.$/yI�bN���?�����)CT-N,�ߵ���.���O�uZK��Fg�p�Ǉ��{N����gj������;?���[_�eF�Ua�rX�+~��u�-s�N%hy���һf�f��j�U�����~��U�%�G�e*��m}E��D�;�j���W (�����q3�����~��oQD�H�`F�C�~�ag\kq�.O�|��v�(�wu�����e���IC��;pI�W�L����ʠl��}�HO�t�ޗ�P�bc;j�P�jޡ5���UJ�}	�e?
J�Q�/=1�i7�'���:Lbр��'���-L�������+G�T���k��V��.x�;\���D9���!e���.n�yG�P|@%�ܰȝN��u�PN y�z�7׈(Gt֥lSIB_���I�SyX�������_u��l�c�?<�!�7x��q��ƻ]ޫp�����+��jޏzb�a^����O֨Te�w0�V�w���l����U˚�� ��f�k��
[g�/���~�B8�#�c��@^T!���'՜/��+{G���~(b���@�M�u_T���QIM���С�SdM7�Q9����@:���ɘ��&�"��,�E���T"��Xϓ��r�UtzV\���o�feQb���vF�7"��S��f�5�;����|u��Kx�t�ֹ�5��V�;�Yh���+��H���&#)r
��=gw����c) ��.�3�~:��
��zD�pKX6�R��y�(��]�֤M��E��n4��T��f
���c�d�P�]~�0wn���c���%?W1�Q�������|õj�K%ր�k��^A�񁀊���5-D�2y�,g�S�k�J2�a��M���C�B<��Vd����HN`�e�<8t��:}�:G��:,FbZt�''gZ[LI��p[6�k����1�Z�3�mT�s602�#%i�pq����<��������g-�੏�zx�8ã۶-1}^6j��Ʉ͸����Fuԃ-I|?{���%6�sƆK��Лf�o숋�o�5bDl��{�"��1Hӛwl�ST��S���P��E�7�\t��}��b)�OW���[���|�Á܆{��Ǹp=5󓇤�d|�:����LPS�O�y�ĭ8�!fA�*�
A�� �V'���(ݭ&�q���P�	��Mx�	�Z{�stǭ�Ex��� g	��*�6Ҫ�a���Cp���a����^����P���?�*����h��N�b��[ Dx��4��MB>��3�;���fvhB/[�R8�(�X,w,@d��d��|��J�g�������bY8�-�~π��Q�q���X|���Y�R�l-�4U��&�Ğ\�ߔ��f�%�bj��4[���0��~��J>����ϓ@�W�!��Y�VV%cV�+�K��W�}C�n��?z�$C��I��c�[�r>A��JF�2�i��a����̲a�,A�C(�T�?	ԙ
�
徑����{��Ʌ3DC��l�K¸Q`q����ah�
������\ u0[�ʶ�S���#��	ՙT:xz%�S'����M~3�R(r�٣u$]�+C&!uο���^���@�h	�����h)2�oaз_�(��yj}#>z�*3'�(�}�Gi��"��&�b�+j��P �M�<��5[�5��]2{�1g7�ԇҲ	�:���[�Y��bG��a*.iu[����F�Ώw0�#�wC�a�$(p�~��V��L�%�u���V�t���3V�{�jM��Ɖ�V�V5vUX>{�W�ѕsQEn���E"�Ԥ��=�� J�1HJ�N���펋h{�H��U�$��9�F���I���Rx:�(�4�t�����tCm2t�i���:�%�Y��{]tC�]���;�o&��y����D�N4a�T��%y,c���ݷ%+�&m!`�gY_?) ���~��#�t�$�"C&�%>굧�>D��ٶIc��M�� �8�m��	��>���E)=Q�$��a�b~�4����8�)\��)��N���@v�	�Hhۼa9e����(A��!���^03�8�zNKsl���:��Q�7v�ə(�P��E��mU���7�����|���Bt!U:�����\h�Q���Y�Gi��xe���&g���`���,g���zV�d�����nxZ5~��]{���(M�x��_M���D���2���uY�
'�<y�йS:����4���SOy��!�&Ҝ������q ��U��w��S^�~m�̦��Bq�V��z������N�~%����?I)��.JW@�̞'�0}����[a���9��p�ZV �tP��>�bl������d�^K;S��*�Х���}kQ�>7��9b����L	���/5�{��8[�V�J�:W](��j�������T�{���v�!�Q�i��e^��q�9h5��v�W�,�x=�W�jK��0���[,y+o0��k!E���9���$x< Ai���"��O˧�)� ��]���}UE���)��.o�ғO_$1��!���*�_/̆ÀdN^�l��A��^A'ƿ�m��	zm�$��q��������15HL�J��C�����"��e[Yp�%���<�T�6#�A�`���ݫ�v�c��#��O���!��`r��O� ��2��$�DУn�\����=��w��,(�fN����0g�xsЪ 郔��O�GWP��Y�$��T�{�T[���p�m���~�4; uD�X�"�3p9i�/�x���1�I���e��V��E6)"��>>��dR�ru@YM]grnQ��!���;&�]n3�.xB���7S<���q��'�5��	
���G5\�tZ���-��`9��̅e#�
��c&���r���}y#p?}�l¤�4<y�=�<x??���|&���2�j�R*��`oe�:k����/t4�����!��I-1��H}�E�#bXM�8��sx�H?��"C��wMJZ��N:axf���0��Ձ��h��v���N����̡4�{�Ko3��>�S���w~ޥ'9�d�0}��~1t{[Yc����0'O	�t;on̖%�s��>�<�\�/�UaV1)^[���D��B�'�\g�S�����cp=�]{/R)��a\^�!�v)+��Mdlx�.`@��,*]w��ҳ�Oj�<�F�r_��1Hˋ����,n���{'�WҚ����X�{���*�bq �	\.ἆ�y*�g�N������6��UQm�e6� ����I�$�(�ӡ�\ǃ�>"'!��`)����>�T�b�:�2@_��)�m�׋=C%o+0���}*��
@� 
ʹ��=.jT��=]��ҽ�.��i�ZJ�,jn��^ެ���*�y���G[a��0ci��yV��%�>�+�L�;!�)y�E&ٛy��Ґ�a?=���r��($?/��8h�,Q�o��\V&�sO<	yƎ�jկ�+�E�e�	7j!'��HZ��u/�~^Ɓ}ݱ�h��O?`�q	nA����5���1�_�Э�s�?��Z�%Ň!����o�����ϯ�Z�N��~���F�U�������G-�؁��X���H���������
r��(�ca�4�n�I���^��~�F�J�.UXD�����E����o��O-1?�BL��F�6�4�ϻ 0n�Ͱ5��Nc����7�������`!��^��@�7�󓮪V����n$SL%�گ��{&v*���� �A�moV�6�7/%qDU��.���j0�lI=׃K�60�|+��ˌ�g��d3��(�A�s)���AT�2܋-sIG �<���H�pk�o�g�+t��S��J�[�	��Ꙅgh��#mM�#AA/Ɵ����(Cg��ߜ�IJ�-kΓ��ρ0hg�Zь��7�]��8���ݱvL]�ҟYNHuL٪�t��N>��.s&�eIP�m߰�rNQ�/]�s`B�����9�;��w����u����-�,����d6�m�N����a�������'"W���8?�^�c���"zд^��ȡ��X��v��Nt*	B��cÐ d�iG���Snza�V�3�_a[ؘ:�vt"i-��7�w�"�9`C�x~�6���D�/TR��S�����ξM�if���Z踚]�w]G���� ҁ��D��R�ՠߎ��
�j	�B5�4�7���6�`��RQx"W឴)�3�j;I�MD�*��8��y>F�T���g��a�2���aX��t6�f�(��"����� ���:e�5�Y��[�N�*��p���ԫ5����z��
D�F!��J���&xL���	ً4��$/��a�S|���{c%���	�"靖/�Xܣ�eXy��'4Ԙ����2l#Ι�����W�g_���%�He�
�(@���Gb����n~���O��Jn ��������3�NS�z��;~��B�>N:�QW@����t�����-��8=T��ֳ�Wy�3�M�A�h�2G�<ޒRYL�����؅�U3+j�m|~��	�D6����S �:7���.�}�D�R� a`�2���������҉�yP*�`��B�,p�2K�_8�
'@���VN����A6 ��ݥl&��&����Y�%�� 6?��sc�)����	���}jY�HI\��*��
�&t���7DQ#��z�!�ǌ��x���0��q�*�������������i
���Hu��0�g��2�i�����`!��b=:�V�[>_�-�Gh��2�5��>�Pu�W;b��2���������Yj-@�y՟��W�:r���3�'֢�
5Dr�i5��&aL��ՋG6�Dy��|����`�R� b���',����mvH��T������6��~O�!W����)]#:���it-C*j�񀐇�������
�� �̤e�$X
��It۠�����C8���)Z��������GԖ�����.I;.9Y���B�Ѝ�3���2 �1a=��k�>�\�p�`��j�����h���t,�)�6�
���Zz��!�1���]����>���gw��H3g�^�yo�2���Ř/��2h�"k0��3i�*����C�@��'�*
��*� 3����8E�"�%�%S�)ʨr��W�Q�b����A0�	av�E�EV7\.G�.	���:0�<�bë�gG��(k����3����c:��h`]�3B�1��ĝ�U��b�]C��VN:Cz�[ۛ�.���V�c�T{����2pK�g�����^k�!�}�xF�F��J2�'j[Nn�ץ:d�3Y��`�Re�A �mr/s�H�0�^M/`S�u;�MH�>��{�ʊ�Y�N����Ќ���j�B=��//�C�&t��;xt	����G���l���BqzP��@�64�$�W!��R`��g�A����[�<�����3��l�: 2�]��Y{p=��3~��:뛐��tDq6�Z�
��+A��Q�"����5=��AP��&� �ͺ�M�0�@�CTrp�W02�(�'ʵ4��b� ΡB�1��a��q9�$�s2��M8G�EQ1<ʐ=�:�uQ�+�]�����\��:ُX�}��`O����z�3���b��\y�f���1���~�E0�=�,6tQ�θ1'2h��n�tZh�~m�BԷvkL��񛆓��a	H���;n�����f�d�-�E���ːo&Z0�y)oqT���'@E��y�՗�Z��� z��Ş6��^��T{$�4�8��i��R��=	��=��+�0��z���"���-�jm��'��zW�'�b���*�p`�p,*8��¶&�y(D���FKHt�����'V+��5����G�S."V[Q��9�D.�rS���o��>>��a�œB���@[�|�ŭ���|�ͼj�(4��m%�S���3팆h�	ن=W�b7.���p��I�kK�_�x�����^�e4<���Z(��:��R�l��C�P�z�"��f
����;F��52UF�:����čn�+͆k{�$b˅��$����=�6�l��B���~Þϭ�]з�YP�-W��8��9������MIVrv���L���g.��f��i/�����t���%us�����@4����YRUjQ�A�^CZ���3K�F��#�b�OA�e^���۴�=���H녫|_c8ձ>��h���d�Jl��1ė���=G�dY�@��gg��A��R�ޥ�P�����}A^���E{  �Z�u�D�f$�}��ě�]����sw|<t�2��s����d:C�d#<��V��+2�S9�2�����C�n[5�J������+_�0��7���Kz�?rǳ�L��v�N*���H�D�c��Ӱ+���F�YD$�T��G��J�qZ����R� C�ձ�;u�m,����J5+��"�Y�zm1�[��u�����-2e�^F��k7z����r�ܔEc�z)��nD��0vp2���q4��~;�g��q+�vG)E���QR0g�/W�2������ja5&��ќq�?+wr�Ѝ���觫��D��io�Heu_Q���H �A��G琵$���r��=��y�l���WD'
�"l&CJߩ]P��$ѓq����VGlA�8�ׅ�i��*�J�4�(FE��#m�a�Rp\z	��0bwB�7��N��3��0 ����~P��� �IR�,f���iui���F��J���7�h]��	�{�N�-���f��k�H���R$v�3I���@�KΒl����;�L��qhZ����.�)Oj����m��U��Y'����t��r>���� �Z��@`�rS�>=A,)Ay! m����)�(�� Xf�J6���n����>U=�:���_�<����gQ��C ^�2��D�-1F���I�,��`��â���{/�N�Y�5>�a4��-�nRb����3Љ2l�P���h�A^%f�uň6�j��&_�����>���H=�q:G ���e?�37x�w�SHw1�g�����Ct?$A��Mx		�m�q魯�-�d�����	G�M�LS����7%�Tg���
��H���E˕���������4�}���Py�)��#|2ȷ|:����.�������>ז��V:�i[S��t�(k��~I{�ք���wK�>|>�M�t!W���8L�2�=�yQ߱Q����>Gj��ag���ަp�;VT]k�ic�l(�1BM���g�c��fA�2��^M�>X֔��x���Мa�nj��>�o��~w>~^s��?����.��/R�M&����gVE��B�p�����z��D�Øz�{��q�D�ĴM�����Q@9�9�7*��?n�UM�ʷ��C��@��_�*�?3Q5 ]!__C�z�iǠ����d<te0��Q6g;���ǹno��]Я����R��3�$6�-�.�z��h,50m��]߭�;�٤��Ye�H=��-�C�|M`eq�ˤ�_���[��-!���E�ޟ=��sPzF�^J��69 �5
�AJ䛝ͤ�`� !M��f�L吉]9��,M��5�u��	Ra�M�j��6e�tN�)�g,I{��������g^�~�;I�vZ��@{HnU.�OR�D���i��!�Hő1Fv�@Y�ش�\��/E�<## ���hY�gTsI{�T+o+��������CP*�o`����M��S��9N������=r��\ۼBn*��5G���$�&�
�r�%<�{�=*i��'�x;� ����ji��A��q���x���rW�˸Pʠ�z��-��	���i4�f���2���=�o�r�Z�r+n3�&t�=�mC�|#��+����b���]�{�˽p� ���6t��%�r�C؝<��mߘ��;�z��O~�
*c������Ƣ�n��2����K-q}i�Tٌ��PH�ŖgĊ|���7T�=Ū0�BQD������Z�\|���u�p#i��*�֧
���ԔAD~�11+}Z�Eh�f�> U��  �Rم��[>e�t&��O�!����?�L���K&�U����=~#�W�ni�%��%�Z7�~�{>	2y�BY�Yxak�ݚ�l,�p�5	���F��`�pd �Cf�����09@�Hb����M�!��d��|R����x�V��8���x��=�ݻ6d�+rI���}5N�`�X�K
�;�Ec�0������u�&�p<�P�2�4rf���vW�s�],�������x�yֆ�v�J���t%�d|��D�;� @�̻�a�M��uv���X A��!��#��/��@���!x�
	�p�}��G��}Q�zۖ�]z�Dw��s���)(Ղ��5	�C�9#	0�0�/�&��xBŠH�a$�z�Ʀ�_p������I������f�Oz@;�!<���1�"��Z��:��-!�>m7�5�נQ����1��WL��4�	Y��Y�#��x�қ�\.W=��6��VM�Ip*�E&yP�e?�(�m��#��Nv_��:ò�u������L&�Es�VQ����5�R��-qU�$��������v}����}�ʣ��]����8��I \�����8G���w
j5PԨףd3K���+2"׹
2IЌD��G�n���_9��p `ggE�Ğ���aT��k^��J����'/���>v�G���V�-V��#��(�������֥�ܰ��d%�>5�i���R��p�tׂ��Asc�3�0 x��{ H�z��|�m5M�{�K�2'I/�����<�HCe��"oΦ�X�5C5��պ\\��0�$o6m����"�ZI"��!3?�2����45+tf��B�-�k��^R�=�a��#����^�(ヱzy��͚�i�ڬf�y Z~��%���Z5ؘ�1G�'�Ƈ����2L��l�+:}%�U�i�J�آ��P���ܰCQ��Jo-Md���ƅ�o	�J�`^q�H �#����B2�2�>�9�-��3���u�"�&�����&���[G5~1eryU��Ʃ��ל�:����TUj��⺌��d6�_�{ܻ�m��A���c���#�E�2~��R�v+�����M��gw���M $F~��"C�NfE������M��Ef�"����ͼ��8ZΈWx5j��3IA����Lk/ש��gEl]D�'���������4�y2]Q�F?��
���GP	 U��\F�R!���,\O��rZ�2+��֗��޸Y"TG\���PT(KS���I`�˯�O����Ab�zW 0(|0�t	�u�ȿߊE|��xZ�rS ���BI��1����5�>�M�/1��J9�P����y$��8�_��*I�5�f���8��yT2�abB3Ùx5d��T'�ҁcRa���db��H�yx�ʧ'�CD���n�O	RQq�X&	��J8=\E�C'`���v����Zh�YS>�	�v��u���M} ��Bx ����J$�%�۵k45�O5bm�r�ݻK�T'z��0D�;�c'c���P�{~��Uٶ��g �V,�xR�|�;�t%L+I��P�ܿ�Jh{�7la�)�B��	m��t�J8s���6����4������H8��u�U�[l�PT�c��x�ES_�Q�E��֗͟�F)�Q����ē00�#8T������Y;%�rZ�9��;�3�`+��-�m�9�ȯ,�"7�Y��n>�KUڡD1Q���Mj�]�lg�M���%3Y�/���6�N˗H�6�~�B"�ɟ��]xJe�,o�_��"퐦��r�=w��������0KO=���"\d����'Z�,F"� �>Z��Y��&̬g�\v�rk} [v�2��k�/��#W��ݼ}8��yW�U�Wb1i�e�� �lv�{�	d�}���b��t��s�V�+����S��3A</�k)�;^W���GY]�}�&�~H�RX];�`#���Y���7�����6㮋9��:��
ڙ6ط�>b�)E�9�����m4 (oj��@U}x@��"*E�r����u���c�+�����^� ���T� ����w���Y�Uf�Y=�@��z.��4�-Ҏ�sC����v�/�5�/ :-��A�Mk��F,�+��%�a
���hN��S���� �����GRR=�M��~	q�-3*�5�P#/>�h���/
�ڰ��Ż_�p��9 �)_~�
�g8?�����#}};g����.��ʹ��B׺����Of�N��c�eM_"%��*<�cyҖcR$�{�0%yX����O>��v��o�9!���TN�kA��qMek��r��'�1�G��l�}H�qSa�쯦����X��D�}}u��?`]��1(���`�r&��\>���)�~u�U��'�k#��*5j���P�[�9gPx��܂�"���KK�|��	M$� �#�l9(���%�[�cC�<�C�V�0l�z�AX�{���1(���ȴ.���EA�u�ł�O�hj��@;&�I.����c��_6�!�*��|�n"����a*��i���-t߯9����.�.�Ϣ��*l�KSH}q�S:.wJ=F�%5n�[��`�sV�Dj��U@]�VY$�cJs���Sm�*�N���s F�SgL:�Qɣۏ�{���e\魞���ډ\ȝ~�3� <%h��<�����rx|G?/���ɇ5)4�g+Q���ԕF7��P3�6֞U�p����D�eLf�gJk�f���O�E"S/���BO���8�劖y7ѥ����Ї�o���Jg�Щ��&���,�_ÉJ%�}�a�0�z�|:�l�-�1�wՆ���]��q��-d��cP"7{��2�B|[M�Gδ�0�7��T������P����-���rR��z�f�*����S5�B�?צ�Y��vLT���UGzÂ���d��+(�Z5d=�9*�K�ǏfxT�mz}�W�2Ɉr. Ji�&���Y�H���>>��(l��&�X-��L�F���b�NzC~�74��C�-u��yxD�fƘ��H֟�*�ԫ�@��6����.�2b�@�ү�n��X�B�d:I~�J)rQ��X�`銘����WpȎ�.�Ey:����$hm�vTV6�O��3�l�g$c���<��}������/̶R�e�"��� ��c����=���b�8�Hg_�S�F��)�?�.�����pt�:�Y	�V���ia��k0h��'�eq�����9�����_�Q�>wӤ+�$�\�q*�x�-�<BJwF��Y�pC,C�D��}��Y���s=zFO��x*0(�x���:�W�F��6��:���S	M&�ho�w%|�R ~��-���Tm0ȇ����/����_�C�|K��%�K
�0��e�⣏c������	�G��ݭ-Fd���!-(�����ci8�im/�0�EB?�P��uo����"���ڴik(\w��W�Ќ��Np�8�lvʣ��cS���uq�]W�d;�b��Fg��#<�=�o�81��c��������B˖�����C%�s�Ao�xyDB`	kp�H1�n[���u�����W���E��Ƶn�j~q1j��^/ͻ�p�����%���xj�~��'��ք��U۵�7mD�R��1�ǀ��j}dƂLH!o
�{���k�;�E@������%]�P�' �A ��\ ׄ�|O�p�&��^�:.�� C/CL��
�z��'�w��~�)],A�Gj�H�L ��}�=�9��1�d�	U��{{qת��B ����6v�85)�_HH����_�+�@������D*/H-QcKA�}Z�Arn��V���e�
y�Ew*��� ��� ^��s�g&ɪ���[Q��/��UTǩ���0o!�MSHZ��M��hlg��T+�}���X�
���e5�jCu�Wa,Db���L�z�f&�U�
��iFه��m���}�I��V����|�$�Z�UajukN�fmC?/_r%
f݀�
pk���
O���ۈ�yg).Ԟ�N�|��wے�P��hu��ElÝ�0�����;���Y�+6	���㶐�I�8,N!��y" � �YG8��-�k*4�z^<�m��A�H��-��0؟Gg.c~�[�y���
1}��5ۭQ�Đ����>;���vDd�q��ze24�Zɐr�a�w�p-��Ԉ>�@���]��~C	�8���ܬȣC���|�MߤS�t7��V�aRh1��Ĥ%���d�Z���/d��6:\�n�[� UZB�a��k���`-�~l���`|�؛�؊k�X��V����30Ў�U������R�	���"�?jc������7"lE�l�����@�hs�P$K�`�1�QNń�����$)��zB/��h����f��g~��]�� j���>�S�q%G}���N�]AFWd
ӯ>f�x��p>ŕ�Yu `L�cѴ>�ʳ����Ŗ���N�����a��֭:���F���B�Nz/������N�[{W��B��M�4 ���y��mx�l��I�#�A]L�� ܆��_f�4��zK.{�|uQ1W�Αu��Ҏ 	mL��٘^��������&�/�<7��ۦ4�=hY�U�����ow)r-ڈ��e�7Y2��[��xȧ�N�����	���m���d��i÷��ӘD����v��]�o���,1���g)����do0���ջИ��$�OO�|��uZ�X�:�pi�ɄTōa�f%��Ӌr��d/'+n���>�P��j_�L�����[��~R���\V.d_δH��<{�L! D�U죅�pLT�������:-�p�T�!��|L!�*U�j3,�W���5�;|��5��7^�=����a�L�Yi�g6��u�ס�m�F�P����ܪ�J򨲐���vn>T���`#�*�40Һ���ģ��]�|^�?�8;�73�|��R�)`f�pz�MM��O������6>N�����y�.s���r�=v�F�SM�P��|��U(Ũ@�p���:�gLp+��STا��`�r��o�bC������A���o�����2uF�7ֳ�%��J$���#�X���9A��~����]��("d��-g:J�Y�H�^��o|��T�_ar���T�_)]%]�<u����w���"I�*��e�3$ǘ*ǟ	����/g3�V`�ir9�`�M��'l���鮹]O:�B��D`;X�
�9X��9���ѾU�,I�P��kϐ��l~q�ƥWw�o����݁��=l�.���M�2�ʒZ|�P'�)��-���U����M�gn2 w�=�����>_�/ V!t�Q�N5СNЀk^:��ۉ��T�o#�z�s7�|�ʓ�n����t��a����2��^o醪�� ~LNcD�67�����_�<�ھk'��57�T�}���l^����EJhF�Rӿ_|05%�����[����h����~fQXa$��eM4���2 v�z`�T+r&H�!�G����ci��VTڲ�q�r[cJ�s�ѻ)���3���I/�@TG�1���B����Q����S�8v�u̞X�҅Zd˟�������o���7mg^�������]�c<��i7V~�	*]�
G��m{3�o/��/��pp���9u�c퍺��4�g�+7}���҄����{��S�­���I[p�%�cҧm2s�my�E?(]�d �_<67�w�Wʈ���C�U���+��]�-�jr=�lGa�Cc�g�'L{,���nl;%���n�'>&>�nQ���V4�=��{N~"�B�:�B�@�ݎ��a�J�l:���]�Wb;��mj��}[��%�X}8lt��j�?\͹�n��z��C*S'nm���&4i�1�[�s-�����b���L��猀�.�n�ǘ=�����x%�Q����8���'��©μ�	�c���iAh�s�E��S���Ķ�7���
5��u`��-��J:����(&�B�l�I�V ���{��J��]��9T�4��k������C<3����!�H+b|�$�,��ъ����@�J֑�#��=��}f�
/2�]f�����F.���Z���"`��oE��l)gf�7+��f��J��A�� D-�%�L9�sL'h_e�Dt�$��} ��|V:��);&���Ŵ�L��\ ��wq�/�Pg͕X|؉^���̢��Mc�W�qvD��W��G'=3[a9�{U��
�ј8(#:@+�:K�U�5B�GM��O�<(����!�s�����_��hB�2c!B�'Ҿ$C��x���ޡ�b��F"8����Q����ϲ�OQd�4�U�X�GŤ�J�*�-�nE�Ȩ��	ѝ!��or� �Z&"�p�~�D��k���,[�":�v�L��Q��k�?�^��CEĽ'l�	�(*oEb���O��w:4E�ѴL������S��Bu���s��ܭ�|�vd�w���l��#��CW{�"[AYC>˪�j`Q�w� ����[Ί�L��k�9kK�`t "Ayܡ����d
�/�͘I�}��?�M�h	h�Y���P��v�`8�!m�����U�OӀ{�֕��<by�PI�ؘ�W"��=�B�<��Һ+�o�^hB�	Uj�R��o���Զ�(uf��,�N���Sq�?6DWΟs-+"r�@/갷�'�o�W$��?����xHZ��!��1'��`%��y~�x�@��9α��i�h������Q�g��_�ⴸ/��\X�Iߜ;ǅk2�u�`���S �^�3�]�o�D�\:�8w�ʞ�p�����ՎԶ�K{���yH�BN��2��"B��]��X���M�`t����93Lv���.����*��T�b&�2��hpu���+$�}�U
��3E�}$� �83r��\t�.��DB���x�0��ɇ4�5��
9u3(����a�	 ���Kã��cy����n���|+�A�|�z4
$�-�bՃ3�8��h��k���B�Ɗ|Es{;�p�AC&<0�͸���j��*�h�]��n���A����=���~����+�� �&�ޢƑ�A<����6�[VO1���ʝ	�TyX�Z�F�~_L!�1�;���sM�:�� {),0��`qNN(�]�������P� P�?�v�ń��e��5݇�b]��T����y�!ҺN�� ��ҷ�KsxL��r�;���`�[rDB�d��I\~��>3L��L�4��Ȩ��q&�Fͦ�,��ݬ_t>sMD���¡��R��CtQ[�Wwa�y��͙q/��ce���ep���@�SV�EXi�r:~΀�M��7\��T���}N`�"RW�G��_J�!�����z��i>R{�[_����o%Kyb�!nc�D;�gU#�V���1s��N�qV�tR������f�Ft�>D�� �Pq���}����� /ykG��`|��.w��lh����E��t��y[�[Y����4��z,�.�,�_�z�u�L��(���W,G_$r�G�Ʌ4�f6��Z�`%��������	��Fs���2�M�H�#j ���,o�g�%���`�u�;t�y��n�Ë+h!�ɝ:�Un��b�z[l�r|�HOS���T�������f�*�vb� @14�Y1��*��b[[���������6��(:��8�Q�!�so��D6��E�>A҆��.��&�|(����P�����It��?l)aq�qnQ��٭2Тty�1�.��6FB�+�i{U�?c��Dy��6�Y�i^V�]�?�t)B���Nl�h���qG䪕����.�������fZZs�q��R�VE�I�3��j
A0և�i�nM0f�Ix�5y��쑤P3ueq��7m�LG@_� _H��ͫ���)��?#v�EH�����j�Ix�qp����xp��z�Ƭp|V�"�$[��h*y��U�:i.�X@(�*�V�2����W�ZZ�B�|r
���DWȗ��nK�n��} �37���G�� ��Ė�$ i%�jV��V���ƶo/.���T����Q}�.��1�{Ns���w�t��n�)��f��1p�?�Y38��ܰ���-�5��Sz��b�D�`"�$��	%uDs����l6��1�p�b	3��%��Z5w��<�.a�xaJ��ue����B`-潘T�j3#
m��䴏T�s��A������Q���ȣ�~��&h#?�2Q#`B�ϟ�'�m�)ΞnB��I���L ��.r�Q��sMsdoԽMe�&0���T��kO�۝�G�T�ff��l.k����b?v%�2�xS8����I+J��̿�ݺ;�� ��f��vF=��bMM�5�c��4�/�D�b��čٷ�x*`��#��С���&Sn6X��9�Қ�Cϒ��}��t�W��~'�� �Z�ٞ]�-�*�S���&�Qa 7�X?�n����w,�s��]7ғޏ�_���
$믂�Ia�<�%��j�A7�6�sMh�b��uп�`�AM+y�c��A#����K�X�b�|�4m�i����=�������j	!��hPݳ�P�n�V���v�2��F��;���nZ�>}r�>�*��Z�@���iHFY#��%��,��a~��vp�DM�,��ҁ���Q���i����V�/�1��/C��=����.qp%�mS�:��
Ey�����\0�KA�Cں䔍֞��-�cӷMw�<�!�!�c�a�^x��<�-�Ĝ�/�>}G\8.2`}�(�蕤
�b!evUt���}��۝Y��v�����l���v��i$�?`5`ZE=A�k��7�s��L�3�]�2+u󒾤ؽ5P����,�>��Bx�����C2�N��0ۗ!50��V~�y#u^����33yk?��g�V�[,X� D0�q�*�v��$�'ۚJ��2�@3k���LZ~/w�-(�Jx����Ʋ��2bgz ��
��	u&�Y������`���Qn\{�=Gb,�	j�uz���2��@�}`�Yꇯ����z-�\4����&��d�],�"��8�7��y@[��n4����U��ln/G��N���VN%O���G�q�ԏ,h��h'�p�Y�<�"�? @�]�2-�ܾ���xS>S�#o7''K��}��<l�'��Tb��9sJ�d�\	F�/["?9�e��;֚o`��8)�\�l��!��I���Cr{��}�b�T�>��xP�[�v;n�T���u[�I۱7��:�/Z�,���:�.�/��Ì%ｓj�Q�m�(>P�MY�簛4�1��I�ZE�&��+ѫs9<���D-n�A��؆�˃FR�܊/�@�&{�@!ڟ��0�U2+Z������Oyi!��cb�pEY�S@/@��=o��2���M�����	�*[Ox6zA����N.��(�=�b�0_�֢zq�#�=	2I	���k�6��f�q@�i�!� #�y���ڨ�A�
j��}Ҧ�*��LՃ�A��&�
��6r�����&����*~�?sK��$�����Kb�}�_����]�%��4i�Y?�v%��;�bCz�k�:����G�N���,�:c�U�:�"J
d`}p�^ܯ�S��څS�:��|^NR�Lly��[���(� �*��m�������m�i��2��f��q���t�R(��5zif�j�
jX� 1�҇�x�� �ߗ'�V�����w�ֲ�_8�*&��U����Gق\��3���������L����I���.���z���7@��������,,�����N�U��v�Q�J�A��������:9&���V�4����U��*�4;��8���RD��M]h��#vBB�`@:̭��&7�.�P�L24�1C(5Å=�M����9#�gO� ��{��fQK��+�n�:�75g�t��;|�{�
ϑ_��RǇ��FG�ȰO���&m/���%}���f�GKC����������ch� ">����R�:"�`3�;[�5���l�^0��܂���wi�y���C�V�\֚�sW��z$�n����ex�%-~�
Y�p�e����c*:͐���q֢i a�F��=�7���;�q����`��I�Q��� M>$�G��v��C���h���o6(?��W��T��iR���D������͆K+�ulq\��99����=jw�KP�ɓ��?p��\��㰊(v} �7�Ivr,��-<�Y������Q)��'��(�xGcV��v���Qry�pA����2���Y�X�q��i6A��������Li�\@ f�M��Z��czƌg�e� �xA�w���)5�P+Z�������3_��zn���5�_�L�0})�E$5�;�$CO�?g0���1������eX(����R�rw�0�!M�?p���)�m��@��K�#�����B49�K9�f\��fw�.Uϕ|�͂�d���A&x[��[��|Q�eи�Ճg��~�����3��*5��!ة���ʰ/�;ECB@�98�%3Kf&��k����Pߏ� ����-��Q��W��@���b�-�O�Q^������J7dh�y�8Nx�u�y.�,@b�$���G3�:�o�, pG8���@0��3K
dVs��|�y�]�Ry:���Mw!C�C�7�肃�iN9x@�P�u�otMi�L\Ĳ+����{4^�!��	�*����vՎ~�d��nA��$ۘ�D�c��5�l��K"ڤ��s��s9��Y�X:���7W�\��� (�GӬ��+�(>�"�G�J���+�?-�����츨'7�(`q|����댆l<���]R��_�qj�>���,7B���JkA�?���n~�cP�}���^����34	39?�)�q��tF���Q��j�����=��cbث�:��|���g>���	d�ő��7iF�1ś�t�`%��O��vPC�|\K������)��[�r�
��C5�rVE��s����jx?��M��V�cd��lIu�Ny����sܾϒmy�ђ�gO&v���Ӓ����pz�?~i7���x9j_[1�t��l�(�K�w&�hvN1U��~�/�$a��j#�N��+�5	����SGo���H�N����ƣ�H������)�cG����c��P��V;�D�l��.%�+D�qQQ�ý&��,����/�?���`kv�f�⩏���ѽ����BG>nq���XI�7��&��'k*jN�������øQ�����8�}�G!�Gη/������R����$1-\���U�p��ϋE-R
�?A Rt���l��V	.YX(�/	2�2G7����]�?��,8i�S�KB��^��&�t��S�%��c8���m��m���mF�ہ��y��='�y *������-�{�/�ZVlʋf��X<�0�@l{�ʾ�{Ġ�R� ��
dP�=b�2Nk�ÂR��-���4�7�ꢜs=6/}��p���yt�F��!�KÌ#��� CV�g���H̜}�/Bv�,��u,��Q ���7�p� x�:��J�ҩzI�	ɟڇ�k�Lz)G�φ��	-"�[��z�O�2�e�Z0U�g�ك?p'C7N�����������9���VQ]��~q��|e(�#�H��� �G�����#j��� D��j����k/c���Y��ʀ�(��4��yL?��	���BIA��(þ�`�J����Qm�OEq{�".��O*�)�T�"ӆ���gb=���[c�n�����c�5�=AVw���w�y�@aQ��-�3m���Fr��l��x�C#s^i���F�ۡ4%T'���h~|��P�6΄aQ­�W�NS@܆��ɐ��/�'�\�ʢ»3�k���~,��k䵍��t����+�D��*���(v�ܖA�-���p�
����\��T��'�ۘ���?�_�cV+�9v�6ϙǓ�Ϥ3c���g%������$`��}�Q�Q �1��S��\o�%>G�5��Oe�oz�É{�|{�
��Cr����E����#Q�a�}B����檯������7����6�VP�	��F�|Pٜ���n��11	����Jng��<�M��;�Tu�}[�IP�6�.c���sş��8vul�e�He����k�[y�ad�u��P���:J�F�V�Jq�V��3(��I6c�<>��)XNR;������vŠ+	��%�"B����ꏑPj��L �o�:���4�����L���J"��}!-|j̣T��@4��x���	S�U����L��?� w�)���I�)���۶�ï �i��?��B!�nwZ�'a�;n���]���<U3�/1B\@3
~�m���n9HP��h7;Iq�IL����J1H�xz�s���G&�÷����+X&]+�f(�K�No1��	VL�^�1kZ@};�1U�S6��8ak���Ԏ8k�����b�F�
��!��,�ƻ�8�7.|8Q���|����<(^���+�Ed����c$M]���xs�	����V�Ju��*�h�l��D��
=I/�'�'a=�܉�h�Qh]L����Q��<5n����+2
r��fmj�];�4Y���?�	ԣ����,Qei|��5҄�k����̯2���yJ���	�n�8I�CW�TRX&d[d��u(��f
���=���
c���7KZ��6���A��'i��/�f/u���� ��D$g�ݔnd ��0����\/f!�^v�z�� \�� �`��G`�B%���+�ˠ��Z!`7���r�U4�chd��^�P���@����j�\\�i�����]N�a�4�J�؉�É&�E>{��^ w c��_g��c_�8��^��U#N�LYU.1R�
b�%t��g#�0��|�Y���8��Af�wf8��d�O�;a�u�˧��3߅aZ/.!�}��!*<�����%�6]���2�F{F�]��D��}4R��3�ܒ�	̀��ykf}bۅ\h��<h ο�w��AJ��]g��S�����oq�?`��)�B��?*��� Sp7�D�z�Ep����.E��4$<�݅s��zC�^P �kMѨ�y$��'�9�Գ�Tt*��ir��o���_�Jks�_��آ��,�-�[0�Η�J�D28N��e�������b�b�VSl-Cn�Fۋ2�`^9~nӾ��b X(�钊�Y�@��o��)k��M=���g�y�d�Y9KP�<Rފ�x��x�jŴ~Q(z �+ݏ�B��=-�O��`�j��I9g�����٢�e>�$7��s�@�g��L�LJ�Y9JA�B��~E`�`��=ғ�"c�2����>�a�X�5�L��ae1x�����
%�ƶ�|Q��U���b�hj�8�xE9�.�	�<|�8�%�Z���q T*+�}~�/'K	����P�/��:���d�p�3�r��$~���VP�J�g�(!)<@��p��Ô�lK��6��竱�X���l@��[7z�4��-�(�O{�U�P��V�	)0�PB��8�AS���e�+��� e҃��tO��k�E8>�[�j��i �D	�x�4f>{��Xz��{ZG�a��<����ݛ&�U�ʒ�b���!y�VXۍ�)Fc���qE:(v�����$�����`0��Ap���ȱ�>�M5L-��-�sj�E2�K�����Nfhp���-��byx�$3F����9\���w�<����5�`��������}XJ������T�$#9j�wVw9��/�`YJ�9Nf�5WcAOoe��+E�ZY�@P)��V�\@F�2�p$�� ���!�4B�X
1���Pc�^�c���,g]�kK"u��N"ҭ$AI4ӓ.�>�G�}����'��5�}�V�����A�I�����#mu�v����:�ךN�{q�Jh�tY�O�m��Ŷ�ۥ�'P�Eu��x�ZL�x�"5���9�u=�'�%��d�f�"���c���@:F��|"kV'9� ��%�\��_*�`#�wN�t<�0��1f�8Sh�g�B+}��*DΈU h��28��bʹ�g��l�k����M��|f?I.�����4�*��H��A=�C��a�j����������&�6��rW����_�ymXƃ��Q`s(�aq'[9 P��ِ�m<D}�9���\��`���S�$�3�$����y�`�e�һ�ƤJ������~.��h����N��{rZC�̖�`D�v���.$�=EJ[=if�$�'6$�Ď��I?w�5�p���_�w[ �)�[,��HO�I^��? ��B��8��'���=�z��L=�����'đ���aj�M\t�^�n�b)V�|�</q��2mYL�@���F΅�uKG���1X��-)�Tv���-!"�-f�7�S �iZCZP���/mY�i��ȼ�[��	g��u���|*7�	�I�}�Y�(�x#nmI�=$�0PpH3"+����{�Z�R��-�㼟g��ɸkS�On��0%�?Y:p�g���`N4�F~gI���ΦM�2�[� ��c��&	��IH�N����oI)�l9�`-w�=��l`	�F�Ƴym��+�='WU�e��xo;*����E��E�C���ċ�[MB%�1x��g�}>a|�J�z�t�
�D3�Q�V�%��e� �G��&���ibۊˁ{�|�g-��JZ�4/�Gݾ����0+���VW�З7��d����Zg��=���;�lLG`!*�|��֧{�C�M�]{{,� �V|}r]b�3m�"��|���peD�w�ה��pz|��W�2=� �L*fvw��mwR�fo�&�l�ߵ_�����X��#�Q��qʟD�@�B�����V�v�}���`�Y�G����*�t��1D�������u_$TA�C`����5
�<J2 `��n-qd��haۈ��:�&O��S�Y�S�.�Z��$��Sϻ:"�����h�li~�c|�=ɹ�V��R`�v`xvO�D�;�z�#�79��}�66�Uzm��m����ს4������ff�%���~_��I��{�/�](���
����!�#�=y�M�U~\$������(����f7_`�r�mṰ��aW>��vrJ�y·�qED#�9y����'����)R���j��Ԡ���x�����a!,�Y�x���	��ẉZ"��|+L�o���f�p3¤R&�I'0�a�3�%+�m
Q�j,^I��d��H�^0��qSꗨ+�7/�}�C)O�J@��0�TO*�.p�!A���8¡',�i텉�Y��GSީ�l��Sb�Uw�.(���g)�qJ-�V� H����A����L�m��ɐ�.<C���@��k
���z������CD��;�ɴ/]���3�/��eH� ��7�?/�L/��R�';ҹ�m)����o;sC�w���D�=�)����F9J��7���K�����ϐ#��1��[p3�^��������G\�������Ӫ��i�ƧDY�-��Uf:.$��?�
����2��dCj(f���*y�
?��\�<}@�!��H���g��y6�y�s
�.1�����F�g^�{k��o*�q"���h�J����GB�4K�z䚀E
�O��L�L:��܂b%��TW�z��=#�O� _�bw1��5Gl�L������W�@�V��v
:��������n�փi���S�� ��CO�2�_�6r���W�I�+B~�����E��б�!]����/���)�.�h���� ��L�9����P��Ɗs�X?�d(�"�/��R��Z��Ϧ��)z��0�Ծ]�hU�'A�Ӭ0�p�r���SDmA�epD����.J[�>A�U�P�����&Z�c�k��Lpf~������"��2^�2s��Û����G�PO�2��2"�N~�9�V��	�K�;T��j2]]wxr�T `�N�J_'TO&��D��PL���'5-�d�����z��B��#Ij�@�j�A?N��5p�G�����]m�Y�(����tG8�{�ƥ�Fw�u�gǾa�}ޔ<^k�c��y�0��~=8k�0�2���v֡Qa�(�t*��+�%��r�:j~��(7c5����cc}ۅQ=��f�"���Ӹ9���d�.b��_H�R���f'ʚ�Ӭ��iř���kԀ=�ߨ]��,�n�)F�P��(��CV��,X&�Lca����+�Ъ��<��k
��s��|���.E��f��.�F���T�ya��_�Ń{�'o[�6�͒�������Vx|Rz���
��~o��-Bc��ʦb1-i'�p��8OZ�f�V�"�_|N�5�ݣ)��������iü[��sbr/��g1��;��aOj�a��+,76�����~ߩ[LPP�Hn����K�Z����i<���$l����]dW�F�_�J��S��9����R�K&�9^�9?����S�-˾lZ��̸�
�<T	՛>J��r4y�~�g	6�w����E4�׏Y<�,�g��E �!��|�Y�����o��u��-��\��n9NQj[
�"����"�������=�x'���%o�3	�^=�l��,PĈ���!�5�qFL�\��f�I�f湶��MSU�!��ˌs�{0Q&�KmG�o�<���ja��E@�G,�6Կ6�w]ь�k斃:��*?Ja뮁"�%eؽR>���sǓ��]���M �q���������v�v1����&4��y��]O�����X�<��?��8ZCѠ�P�5�)M1DOڄ$$�� ]�^�Z���Ē1��J_����<�����t�L��*��&��zU���$���1��ߔ)�R�|�yӮ�xo�}U��D�]���Q]\-�-�#Q:XC"� �f�>T���w�3S��9�KFU��f�v�{9UQY��^����-{8"ۘ��3���
?E�����-�fQ6^��쥾k}��F�K�^�٢�s�{#�26��B�i�� ���Ӥٶ�Iޟ�B�	�β��w�z�8�װ�$�[��u2�+�بX�4:}��0��x�ԍq�6�2}8\j/)̣��	����XgRPY(�E�K��#�{>���Pp"�4�*D{aZ�����$ ��5�]R	��G�L�>�!��:�E�I�,�~�� ��u#�_H�$#^�?��f����2��m|����D�n���^b��g?ަ�Hx��]��J��8��,l�K��M����ߴ�%n�H>Mz��UM�/"�䉩7����BN�O�Fc�Jn�\P�h:�u���]D)�8��X��@p�/�~V���xLg��q�}ۊZ�,��CZݜ��֪��n��1��K	< 6��ek�j��T�����b�oI����Z�$���5�N�_�ȏ�y�9�xn�FP(��b�4_)��ȿf3�vbS�����6��aV��	`a��ا�E	>�t>l٘��J��m������~��z�m����߳�.��]F#%�r+NVlA��b ~"�"�y&���0�����0�|`.�+F<�l�Y�X'�ګO<�qHc$A�M�12g�O*���fe����J[�ߟxg2}J�"��R�?���	����Jh>�S��=��S&�����.� �O�����q:b�R�2t���kj��ɀ���sK��#|DA��-��nɹ�qfLh/JJ"�%�8���=|n���$�.:�q�G���h�4$^iiޜĳU�g�<(�����_�@{3V�#������>H#��vZJx1sx0�5�N	V�����0*��<!� ��A��r�|ĵ�f��A�󤵭)�ǋ���0�`�8|��o��Vq�q	Ӟ��U7�J�hg��a]�z.1�a�4HCpJ$W��a���M��?� IS؀:�v"��3���߳a��:���r@#i�˲&��e�8И@a�2��6X�����@���q�r��\�'����wŉ͚e�A��!�ؿ��i�z:߰�����0���g��!a���G�TW�<��-���;%��;y�ē�z�v��G��d7�����k�E�%U��B'>�d�x�pu��v)��o���d��+G�{䩈v��Y��.�t�ܓ�ĩ�Y��	��*�ȡ5�� �KAJ0@`F>�-�	-�@�^�@�6c�P�B����|U�����&��=����b�����C�~�f�E�m,5�q4t�����vU=�r�?M��V�J�ew���v���0=jAQ�<��������=��sU�M=_�D������Y���4څ�����)��2mٲ�o��͌�t��(�5�Wp���5�)*���((�5�;r[�A7_ �8�!x����/,�'�:F�<��������P*�=���x�u��T0�d��a{����o�y�����%*������vXb˒KE��[u�Na���9�^ /�����_Fק � �{�%��y������830��������+�)�~]b�4䑨ŀM�.��69f:~�If�N@{�iGF}�"���)��<q|q�894C<a4�I���b��ӂ �g�Z��%�CZ�<s{�pCw��:�fCہ^P�:db���#�8t�X��$kIhH�Ȳڄ+�Xf���ٙ�T�Ŝ����.4���ږC�m�A���\epHhb��m���j��cx�	ZX�_�6��7����Ă��5ٕ*�Y��ik�m� $Z�����^�c����-�JY���e���)2(���K�^�l) �f�ш*�����g�c��c�5�b2���dK��%��4�~���H���~��A֨����(��2V�#{����e�H�6Kr^I��u&u����b�n1��fw����h�+,Imz�^�Bs_������|Lpȕ�EB@�����ξ��40�g����{,h��S�6���ɴ���O�֋�Z�~b6mx���7w���!U6ԜC.V=�c��We)�|[��H8g��?]R+�e�������J
�D@ǂ��&,>�����u|3y�99�Da8jc��~#%���{�x �u�Qj��Y��*�yk9�L�?�E�Uo��:Gy�v��8p��fZ~���j� q#Ap?�쮤�s�ء�͘�ۙ�W�VE�6&��c_9Cc������~�v�rԁ��w�oS�0�z]�=�"��0�㡱��]���{��6�|�ߢتx�OT��|&(>D��Q�P�
Qo����8�85
�n�	P�i!dN��Y59R�7j;"�&^A�|�o�X7E�J�����:�zt�Fc	^d*K��>O�+l�҈���V=1!02�u� �y$�}a&��cԢ���J�����Nߤ���2�C��׸���[�(##	q߇��5��}2�9$�D#�K�nT�ȷ����h�0nK&��ȫ����v��"�K����Ӓ��{pH��g��vr<7��'��υ�2�tO���}?yD�.���d�(���ld�^����O(��_�X}�����������q\��R]�ZH�~���4��{�2���H)὏������6D.��G�,�,\�؟t`�@e�� z�r��tm:��O��G�6�IRe����}IS����M����DW���F�ҳ��O*U�
�)�`��y9ON��= �YD��Z�D.��FDE@M�� �F�*v~�۠Ռ|�]�D�^�<Yù�%��Y�����0��#�"Pk�_>���3A������d��)R��s�x岅 �0� I�6���^@�A1����G%|+P^}P�����m��Yz�-栖u�z����q�eJ=�p��,&��ߚ���?5psZDY�J���Q8RQ����pUD]�y����-�8��#ޛ,P'�ib��FS�cX٠�9A>��\�c�8���ʠ��)z�P�z�
!�i{ɹmwe���L�M�����F�Ș�Ml�緜h?���4@����_8Y����!ϵ/�4��Pl��8�%h.�D���h�3�ЯMw��r|�r818�|����cF�W&wB J���+�[�jm�q̑���V��d��'�-�LS�um���MΚ>�saHo�8��{�F���
T!���16�}r����t�Lt���֬#�U~�pO�rjr�&=�
����*%�?����Z�)?��5�/��e.R�ȽI�y2��[Ɛ��ٿ9�QHWq2���SF����Qg֏�|"��"}N��ny�Zm��6�&�����d��u�"����ܺ{r�V��a�`��r7��J���2n\������q�9������]ma��17~��������ɻ�h�Ti�������-�b��'Y�"W�4���n:H����iC�h��i�Xa��Ua��;�Rݏ�2����/-���1Rs��1�˚��V��L)���f�c4����kf<��0�`���[ږ�;��Щ=��lt6�&�����͜�\�ux���9Z0VH�|׫��[�Ynu��b�����K2�(�d̜�����"��s��\n���1f�]��B�<�#���U��p��)"A�����,��ޡۡx-��	��KKM�=�r�8��Dؕ�A�wKhU`Z*#�Yۃ����R�TW�=��[��#�kE9�it�E�����AX�036�߾Ȃ�\�K΀k�n�?^!�uVA��˝7a��=|��$D��Ģ�x���i6��x���;LB�� x8��g�S�Ek����N�-\����3aR��,���߹�}e�s�]�$�/�p�I��4A/�%�B�#͕&�b�mGVؗ���fD���'Ch�:ie��`���DuhLS���{0z��W"�S�D�@ egʟ!����#�5fDrH_�}��Bb\ :8I �*�?���Ԟ7��x��	���Rz�h��vC���(��Py���ޟ��� ~�KF�M�-o�-�Q�S	l��F�@lk����1�֬EVm#��{8*�N��R��[x���M�}X��ϙ�Z�������:c8�1N\�����:K<1�N/�B\l5�|��x��u;�=��<<���۲��0���V����� l"D��z���&?�Q��p��/�@�V�5u�Q����3P������s�u=|z���Y3�f�@�v>ӳ0��Y}���5d��hg�oظ�D'x�2�Cc~Ϩ#|�5������Z�5k �\����.�=�1���j�}�W=G���[Dv�iQ_��m�Ք=�����sZFX���-!:yQ�vU���r��-������=� f�j��T]�|I��ɩq/������Nbl� D�k�|�U��R��{���2E��5�^L��ʖY��=�_穩��'��=j���B��;�^N8�y�Q[���dk���q.A@��&�������z�?0I�ݮZk#$�>����R��j!3ʹ�ѓpR����Z,==72��J��P�5JR�t��R����b^��bu̮`xI�
O�� q��
-�r�����Ց�C���/Ĉp�7�$���hR�X�7�F�&_f�/�������J�݆�2�v{<��!$Q� .(��Y8(cE�:����C�e�m�ف���6i�>LY�\E��߃�����]�=G�&]m�PK�deRs�c�z�2#~˦���xĐ�#t|�-�#A�"`%9�.��������v���g-,�3wS@�pB���X�C��p}��k��C�Ҷ�hSR���,��ggV;?�R諲Q�e��Vcżo���i�r�s�s���^�?���X���k˳��4�3��w�0���E�V��:��ԗ4{�q���T�5��ર4�`�(8��ֲb�O*�D�7�.�T�T2s�N-�k��7[�<����d_D
i�.��_ �M��UxBë�)8>����X�q|�u���V��咻]WU�QJ��N�!�x�����",(M�4���	-V�X�|S�,��jLb����?#��|�*��NcY ��U�wU ���n$�����]<I�n'��晍�X�=��*uA��Ұ�Jc:*#@b���2`b2GMgmgB$n�~X)DzQW��B]��sd�0z7�k\I>A�6����2�C�����x�kh��kB"%��#'j=��.1�_:'B}�[�
`�/\�J��5��lc,1�k\f�͑��5Ql6��G�ں9*A�U���X�f��,92T&�/�hD�oq���|���s��o��,�"��� h��X��$]�!|�m��	_1��:Lѱ�-�U�8/�Hv�>(+�29�����r߂1f������w��)p]��=�&E��{Dʩ�	���ίC)\ݢQ��>�:/���N�c�
V+Z�$S*�W��>�(�;�j?���w�$2�*��CȦ$��<&��Ou��]��2N��{0�|�������;f�]8a刚w=tj�� �0Uy0[��s��N�!��g���k�{���O�Q�Yv�������(0�VH��|D��Ա�"hUƴ�� &��+��+�lO�Ǆ ���|C"⳱t��WV��}��� �?S���"���(Y����p�[�fQ-��|o�������l�7���0	��q���G� @R,�YWiu"f��+�d*�],�Lv~P CBs.���Av��_��M��.��|Ļ�0�ϵ��e�WG�����2&?�]�0L��$�
�on�<�����f�X��4��mW��ǣ�C��S�f(�/�_�f#	���5�-F<n�>i�9a�)\P!z�+���i4o���$�'}�M6/����%���6�D4~'���w�\=�(`��-�[ܩN��0zu�CF@*�*�k��앖F5)��d�KS���'d�������?����▙]�R�W���{����UL�c�=~��!v��=\ �gOT5���jGJ���^=��̪�Q�yI����hٳH�]?�X8r�8�#���P_��Hh	P5v�:����u8I!���W��+\�/٦QQ�OcP��e��U$��Cץn_��w3��g�6���HL]���B_�ͭߖ1��¬V���Vy���HN�����칉Ŏ���DR��gp��>c��[�=�5���TgW�!,��i����Kj��
yK�4Sh�\���35���G��݄>��Rsi���+[�MȜ�Z�^gn�R^��>:�_s�D���6n?��[���'�OQ/�S�����{�2	L�|+�ވ��n{� Uc�ʞX/�{f��4��vx����(��W�}>H�
�
�`0��Bxu��o��>~��A|�Qh�:��F��0��G�����@M3����r�B�jdGUa�דPo� nHk���֒`��ɤ���}�(R��j�j����z��D*�����j��/��݈�<q�NN8�,%�j�*9��~ڬ(7�y�>�N\�  p���\*�`ͺ�w'�?�29�2���FV�h�V@��Ń9��_E36�V���*��M�+&T�Bk-N�{�XT�'��HO����39}��_8ѕ����`��	���Cy����X�\��M!��n9
Frn;53I��)'�!~}	zÀ��5�O�i6���yȷo�����,�W�i��W�|�M �bA�.��UT2�@�_��K/X/��������E�_�����p9�ϰ���KW�ɭ��,!�}aCJ�v+�H5�A<u"z��1~w�^���.ē�����Y��Nd p�=���:��Ll��&�dk�J�O�e n�|v2���8�Kv`�b=2q-+>z�r���j�6x�!0�
�˩�`Z��aʶ<]n����1�n��F�7�3�}�V=��d��J=C�7P#�|:*�3H1���uY�¼p����O@����(��5�8I�C�P�]��B�BrU/�N�(�K ��<��gnBcO�J��(��3̋)��C�b�ˋs��92�-���y�s�Y��&U���U�6n7b��1�	)t�J{MUG���֟P.���
(Tw�p�|`���,��7�kz��0�T|E�V�ׯ�.��{��>���I�|��h���CfH���<�Ɯ*��&�A�:�C��d�u�t�I�� `�O�����n��6ОCi��i�(I����ў\��K�ZY"z�K.�\G>%���0��F�Y�'�J|L��׮8T���0dZ����D���ac�U�(g8f��.sV���uH��pNz@>E\��QJ���υ��'�����B
���P3��4�|����ƨ�7�#��j�7�4}�Sp�_l�*��n��C��2ꌝiRz~�9�=��;�.���F�9�cv��"K�g�v����GT�6� ���iXe��"��KI=L4�� z_�-���p�|j���k�JW�}�a��F7��\��)����#eh��5����'��L�ܡ4�Zۜ%�d���t���Ȧ���Q�y���PY9����g:\�j.����PM2�o�s`���}%_�[���j���.��pM�F���
�Ji����+�9���a�-qI\���T����\�K�ҡ�	p;�a����T���SI�bX"X-���ؿ�d�6�������3��� !�����{,ٶQ�u��C���с������!_�z	�7�؆͋��.���6	Q�n#W�!7�� �9 !ݯi� c!r�=��%d�/�E�>R�k��}U�q�Ƥ��A��4�Z�3s�YX�;���o��)aoЍ�4Y�����\�n�W���F���@[�M�r�g�6�(]��|-��X�#�����l��=����}�Lǋ�Ȝ�j����k��5N]T�Q�/����%'��C1�ɫ�	Z�3dx�+��c��>���������G6����s�4g�o���y�4"�.Iy,��W����u��6.
�J8��-PA0TW��@����S��L���b����p10��`�+�vg���Sh�7���iB/���_���H����r"9#^|�c̏�½bM�<������0�V�C8��>e ��M�H�����5_8C��+J�1lt[�ٱ������8|��W��.ޟ�	`�p�1D���ז����B��T��@�d�S1۩7�_�<B~��n�~r@|E�[�(�m��S�#�,]��u.h�b,�X��Q5��1��0ԣK�q�Ѩb2ǰ�a��v��?(���r<�T��恝#�,=Cr����
ɫY�x�_�kS;���a9�+��u�Ixt�'M�%<mqq��(���R�b�YL�C�U��<R� ۝uF����Ib��v��T]!�y!��Kw������?�9&� B>������wvwBu�uy�h��?��Z�?�v�B��W�ҎK��4ts�F�
z�$�ئD*C�%��@�a��+u�% BG*�����B ��4�"��.�/���]
-KL��Z��m
v�����F��'p&@IM� �	������A�/s�e�Q�`V��y��Ş��%�m(�Z�;�h�i_������(F�J���̧�ː����̔Ğj��4�ٌ�nﾥ�IT�7$���bd��`���\���X:u��Dm�����B�:,>��C����/���F��$�͈��vEJ?�l�.h���#)��VHg��yZ���M�dy�ȅA̢N�X��03�	�3_wŉ��I:�Q�6�����^��Y��-1�R��4c��-�}�43Ͻs]f�5�	ܓ�9HF�B�6������sU�;n�:�fz���϶�s��"|&ܠ8�][��#��z�?\)?G���0gß��[N�N�j@�����B�ݝa�f�w��(��_�a�������Fd�l���i��� )v
b2c9B�^(��Dv�$�Ǡ�tJp�Hb)�k�dJ:� �+�:��/gw�cS��{��	�\�T���(�'�;��x�\	�ʴa��͐;"��\!/8�J�P���A���kh�j?er�t��1���<�UtQ�*�!&c��w��˴7�(@�sr�����b���*�&K�2h*P�ś�Gs7�@�I	�5���-��ӂ�
�2z�i��R.�Rj���0w��r�A%��v;���
+��e��^|�[�; �=����P:\�[��@��[�x*�����a��*:�@�c�v��t��Q��ޡ܌�A���U�o�
��m;=���i�=b��)�MmgG�l�jy�B3�(��Or���O�N����1:�@|tn	`P�9>�}���S˚�w�n��)���cè6��Y(�0�Ds��K`A��WɁ`����bV���d�,<��9��-P�DX�1��̖�pm!1xY��F������J���))XN�$�ї�/�4��!�6#qD=�O�%��a�̣�2��KJ7C�a��Խ)=��n2p��߶ V���r�̃�g(�����;����#E+kR~T�0ݳe����1��ε��V����70D����,�i=;L�I�%�n��4>}��p�w���^�K�В�K�I�@�o�N?[[��2�T��/��c�u:�W;-e�#�&r�o>���"�s����=�$�J|ba���؉p����W�j�T�s/v�V�[�8� y��ڎox������HT�_Lj�ef�e1�z+���u���2o��s��ʨp!>��Vʇ�?߃����gV/�㊳k.=��.#uKXDD���7�H��g "���{X���^�A���r�raZx��@C�ڲP�����E���<�3(���_����5ąX�ha~.[�~gDjF����C�Jd �˧{��@'�aE9h���TB��NU�ʰ��oC?q����aA���$q �:zB�w�b�3m��N�=W{Ѷ���j�g,&N��Y�;?P&0HD�Xb[�pM�
�l{5�!'�:[.Ӧ9�t��J�������逧S(Q���3ş��	$aHp�^��������]��'섚����|L�v�|*��@��a�sG�l����J38߲-���Kb�}jU;��_Gj�*��6����,��:w?�[rp��kG�(d�:��I�>�}�
��p%L��&艗�r�lU�K-�Y2�Uʝ�e����tHt�+t뮅q�����J���(Lq��:�ɝ\��/#6ʹ|��(��bY�����G�L��lr�X21lyt`���I�#���YJ����Q�އ�̋��uA����7б�!?���H��A���jUOVX�������P�N�`C8&�6Kt�Z��� a��cPN�ѿ"h�=�-]t�#N?s�����|!.6���^$���@u���=�}�*:�bM	I/�f!���Ͼ�Q�og�IM�X�fD��t�Z�ﳃ\��i.y��J���4�����G}����O���^-��)g�{���r)�%ёM�[~]ϵ�(����f���a��O�<�գ�
3%7Ĭ�����'�=t���/��n��`���B�jI�beA�D�àQ����`���h�WQ���)�	���F���M2���M�����:r����kI����r����J���ɍ��>k)���`1,l����K
�5�;B'x��"�	(�+�\b�)
�csp���������Ԕ�z�b>��;���(�����Ј��=��>XĿk]��U�v:#��~���{pHa�k�tݎE�'@����hF���|7Ǿ�z�dP�rFUq��[l�ft9�Y���z��Q}jrf΂�(��fO�[O�H��ubG2�!�O,0q�>5Q�FkN�|�\�ݟ5���ק�/��$���$�q'�����i�7O۴/�в�L{�R9	���#�ɨ����N���m�b��``1���ѱ�N>y��׫��녪f�͒��̀�8����K��6[-�hG{乬�Oq����}ZF9���/ǒf�i�C���E�$�	A^f-v�`�|�l{7��(׵��"~�;���i��<>�,�ʺ�ow)��Z +A��N��L��p��ȧ��in��Z7�+Y:�d\�����L�c���6������I�}C��Ir�T@��_�p>�c6��|B�s��� 9�m��P����2[��ձ��<��@�C��6�ʍFd�g��o?ʰ��×e�<�Ī�j�߄�d[P����K��
���
���4T��-�=�_�^=�C�o����)qJ6��Y=x�ؼ������+;��5�(�K&��;ޓ���Kp���$w�#T9�M���o� q�9�۸���i�Q�)��e��otz� ۋH$�A�%��ʁ�!D��`�� �->(��]We&$�aP�ˏ��޵�h����`B3H�4��ko�yd��������S��7F����sǵ� ��	Q��#�5�R��� Ԣ,sD^�P%�We��u*�<���]�_�sr.�i���i�)�#�#�-�O�����O����8�iY1wY�8գ�0Q��N��?��Vm_��(��:o.7
R�3d�{]o�G�|n��E�� �JS����
w�#g.���'��Ξ �Wp��^T��0"Y<;p"�v�h��\�~�I����������[�_����~\^&�<�1�6�"�0,Z�����jaf�x���}��j�Zb1�:u�>K��B�(2Ȅ��z,���2N�x?�g�:E�V0�j'a�����S���i�<<1�w�q�R_��+S����ƀ˧�˵�t�w_"������YɥO��������*�֑���%&�<����k �U͒Ԝ�����w#���m��ū&�z)*	�p�rC�m��<5�&^<zӟ��/��J2�{^���5ǇšX�v#ut�
,z�{+�[�5��>��\.$�-����\i x���+�I�Y����l"����
����:���CM��%o)��~4Z��N"�Y�� JU1;���*��1~'X����Og�ƍ�D�6&�sn$֝ό�����j��,i���D��\߂��GEo����{>B,��=h�;#� pH�)_��cX�M�dQ��BVS�n��Hb����S�,�϶�M�+�l�Gʃ`C����붆k�r*��%���H℁�D΂7��#_�t%9������w�qm*	4�[�N*�0��E��W�8��C�V�B���T���v}޳Y��-g9�e�ckOo^T�!Bj�_r�!�o���{����iv�6��*wz��P�&J�s`�i��,7{S�y���n3�,�
�7�t�����.����v˸Jh	[��!�G�O8��d�1w����B&#Xz����yK�\���p�"�i���g�]�V��C�P R��`	ge 7�b�LO�{��Γ�YQX��Z[��Z�
z�_''h������2�i9��N)�I	U����g2$�J��/2�:��N�9n3I�(C3;a�L�j�s�*卙���+��F��r����G��;@��'�UrE.���.p��)�;'X���<�%�A)2���E��|_,��µ���L�	1b)d�Fz�����宠iW@�C�!;��� F�ң�f�l��K2������*�Q���Tj�2t%��\ew�*�k%�a�"߁��CB�,N�m@	���;��<K7�G�7A� ���O,E����  Ͽe��zT���鄲@�o�%�v]��#]/��K�J���M�xp���OY���pɞ2�*��91��Գ^�>?-�+e@�B1���fsx�]W�������1B�4�Q��|�4��m����<�����M�@�[���W�n��?"��f�%�߭��I.�3r���_ɏk=��{�W���64�n��V��
��m�x|_��� *!*�a��i��A�.A�D�2�,}�9�y�Sȅ����*|��q�:
Uf�0'�oM��� �~/�ʨ�eE�����O�����|a���E���\�V�Ծ�'�f�,­<�_��&�O�Y2(�@e��x��/�����}���>o�$��']���� ���S�_+Jõ�s�;�%!�����A�f0�ݦ����f�K��!������p�24�F*	��h�d{|*��o�[���CJ��=�=�n?`h,�iD/���/�{����wUy=e��H�SZ�Q-@�\_Bv�R���By�1��C���ql�"򕪵���N30�����֯$I����p�P�B�����Ѩ �����ӈ�����m��j�(�R!$��Q���Om)t�'�w�t�U�[�r	�{H�џ�6��;�U5�	g�P�v�6�_�#70�(f|����%xf���_@Q����.�~ZS��C2C��M�s����9V= ��]�4��䝫���B6].G�3�.2!*�[�nE��2)�S���WK����"� �5�4^��4��S���F�!�'A6�!�|�Z ���,a�]/n|�<������.Ͳ��}��P��&�'�ef=����v�(|�3����1H��e�k��9�c�C�uxr$<P�W��hRa4�����6Q�9	Y4AA�cd�=�B�F�Y8�����P��������M� 6V�"���t��"��4��R]�oh�p�Ue��-5~v�l/#��\+��^�������#y�k�߂t>e�P�~���#ADV*�x����ɀ�(̀L���@U9н���+\�mJ�uʡ�kd� �H��ι 1.����B��7mT��ug��[��+��R�:w
#�F2N`h��qML���w�#�\�Zb�ed�-u�z3	HO��1W�����
���_�[#�.��%#�c����D�O���I�]��n�@���;9�Y��L�WrO�I�����ap��7���/e!�R�oK����5�:� <k����k� 4cQ�5#��.�>��}/`�ݟ���\9	���(�G��F�`���"Tg�g�QyJS��B�4UP�Ϸh��>>u%��5/�;Hh�B��O_��e u�r��lm��T�+�Z��W̤V�L����ox�Ͳ^f�H9	��G����n#ȣ���"�v@�����RNX_oN&ک�Id�����)���~���U㋬��<�K�Okh{��E�����^T�]���/�ߪw@u?�I�ԍI������~'�e5�ƍuV�FPں.cÌe̊s@jcڋh�Tt���7Ӈ7	Hk��k�'����|,T��[s��="Z��گ��V�\�C��?�G�I�Ft��s��$,_�3	0��B���N32��rA4K�����OoT	l���:���e)F,��U�i>[D�1k�ʹ��{EG9��31���v��
4ƻ9	[��d]My�m�t�ϔz��|.��'�P�":N�}[P#y_����"����J���r�y^e��!�"�Ӊ�gY��g+r�W�'R���-ǢS�Ӥ����H�D#y�K���c9ҙo����;9^b��t)��w��F�A��r ��t�P�\���!hH��)�:�� �T��1�v�^�<�T��BG�]H��I҆�);��f���,���p�trY����zל�D�Tk���{;k`���3�`�ߵ�|��L�d\���Ƿ ���(j�h
��怋
B�6' �r��"Vk��� ş
�&)#R΢�d���Q�7�2���:��B�#Df쯊��y���Ƙ81���V�{��tR�i�"�������S{�n��x=V ��2ar4Wӌ�%>���q�;�'�^��h�m�_0������y��x�r��z�J��6��f�t���A��x8�ER߽G��ץ/��D�/j��/̑b}P�g�~�h��n��L�?������c/.�A�(2���V*����ȓ�����P�Q�PBhT\��cݍ��+Z[�j���	��Qɡs�C�eǶj�s�w��'K��.�F��ǋ.�d;�-٢��MH>�崎�Z�B���	��}K�wb	��I	��G���i�(_�sa
��3��F�n^����k��H�ɂ����s>��
����cm'F`췉�0�1�V�	���������=�.����r��|�����ov-Ub��k���Q�!���=ܩ�Q�-T�6QN?���D������F�c�jv�r�6A?&�<	�]3&*נd�f�-k�����i���n��tc����QbW��p�iU��(*=��t�$���;�,َ%��~G��I�R).J�ZO`6�Ǆ~���f��И����3�ȁZ�#	"�Z�e�P��y�'5cF�6�E��"�>1��nO}���#�øv�SǃaV0�4��2U��2�2�A"�]<j;`ݏ}ƕT_M��|��f��[��74
�)5i���3��L���{^�=~V��{�L;���t��=qiOcK\t�[t<��ׇ� ��,8{�;�a2�쮇�N��ZQ|��E��G��������C�_B�! 2�,����.~6��8�bDlF�g�t:Gr���9ݿFCS8����\��Y>������x�Mx���p!�.���r�s����u������t߷8�+��X������?�g�&���Ll������6�5�\�ï��I��
j{������j4Ns�=��Li���L&��]�iH ��3iнAv���U��D�_�2x���*#L��j���&�e{�gf�I8g���������i)���r[��o�)�K rޚ�[w���!�����!mY/7�Ș�<��G	c�Ap��ĉ�h����p�5�8.$�:U�2f���N�F)���۴o���'8T���)�Y����M8[�����l�$jd�� �Z�j���vU"�I!Ć]���㓩Ǹ�Q�PS_�Q������1p����V~�Ƶ���E޹X7
�d��g��[G�=�g-T�&"�_�&�m��\g�\�dː�ƈLʩ���x'v���g�/�8l@R&��5���l�3�Q�:C�t�y.��p��+�C��9Px2���E���Z������#��˙��t��jzc@Z�Z�ӭ[|��CrIM�}h�%B�|G`#Avo�}��r�@ϸ0)�lD�"�8���B�I��UЏKh�;?i�օ�q,�ig�w5�v��\�n� F�Pv&Р�(`)��,�d��gn�o��~�O\m^��
��$���L�pOFW���r/vLω�I:�=L����:r��{��\��oe��L�߻r��2�=?�O6p��T?K��E�뤄����U�
��=Bl�p}�gS+e���� z��[��e$r��$��yT�-�?���ͪ�^�#�U�*�̙������Y*a��m�����l��ܛ<߅~�}�2�&��׭�'��ޣ�g�J�p�1�5�IE+k�a���$�{��D��B�-��E�5�֐�SC}��U"�aa�7�W@��y^ه��Ő���*�1.�����y�D`y���9���G.*����	�%���m��za��{��e������sN�e>�A?r���"Ek�<�������Ᾱ5�������ޤ#G��&e'S�Hu�~��̗�Q��������/3�׀���;��N0�(H�f�~�	/� X���[����� Wu蜃[3'[��������
�ʠi�rD�$^����Uӣ�?�d�#x;`�H���d���,��{�� w~ ,������~�|nMkͶ^UTR��j�����/"u��D����0J�q-��iw�k���6ňF$���p;�m�H�������SD�⾐ح���+�ƈ�x�;�1�)s�ʄGf[�@9	��3X��%������P�)��k�zē^V"����<ب�]���4k�J���I���\�X�HdT�'�12��=1Y_��!B�IG7h'��zIf���]Xm�-^߷B���ͬ��m�f ˬ47��&�n�A�di���\�W�?���L�	���Ts�6Ŝ���bw�hr��<Xq�U\��ߙ���!4�?޻l�BG���YԊ�m��/���ǝ��_K"p�(�K5������]����ǘ��.���/�B�GЭ£
}�(=WL?��[��2LG��X�`[���̈�ГQ�#�N-�-��}����A�R��~��a�^@��g��o�lj}�� ~EY���q+����H��0(���~�)lH{�H�z���_�9��@�}م�ʟ���{s��$ˮB�E'_~v[sS�NRosE�	���8tވ;�P_�sƴ�eӴ�{�*q��4��'��v��.��X��lB9:|���`1S����R�V�?�-]�2ʇSD��i\��V�y�{�ԃ��q���(��&*�PQ�Z=!�>��p*`�a>���80k>3�r���qK# �	U��I�0�x˳�Z��"��u��#��=p/v1A���(��xD��1����xm�����ib$���sm���Q��+��d|t2��
��v��qdF.�R����J{�k޼BMߟ.v)�j��F���� e�Ib�9����S�5��^��{690�
\�$�v�)�ja2�AV�S�bF���]˰������Ưl-[v���O����}�:p@��V�����a�2�J��ح���6��v�v]+��.�m9��*�O�L�2#J�=_܌�!\
�nqZ8�����ƫ��R�TA��5��?Ճ=|�� ~���.��sa5�5����2�
�������ʢ�jO��{�8�Q����mx`�Rf<s�����؈��ii�O�EO�%�m ���B�5��(+�~�v��~�sD�!����B��Ǒ>{�\u�b�̅�wx�N�@��3�H���@=&�H�y'���b�~=!���r�gx���B	Ϧ�ЁSz��g�۩�?'���w��!��P������ ���4jzfB}�M������U��f9�P�@��(�����~���O?�tLBCl Cݒ��x/�u�$��9"h�`O�8��q�T�<B����}��oB���߫�U_��_= ������C_����Dbր�ݖ950���D��hʖ5��(����~��1�s�	_����(�:%?�a<�rT�F��M'dj�)���;�����*lhV�c�/	S��r��ª���]m�K7d�s0�qg
���_���.vw���D�r��'�	��uEB�/5y߉r7a�)�"H��f�0Kb?���X ۪PŚKXã>k4�)�%G���ZNd,�O��� w��������}��*���Q�'��N@O8+pQ�˕�4?���'P��n{�����֜��-!�"x����X�u��q̟	� ȼ,
��v��.�/�3�l_�������[�c+�-y���~#�F��V���b��
/璅���� �)t����u{/�~�͖n����2���GᥛR���t�C�V�0��5S�zO��WEn߂�.�䨶÷��13�W
��W���&�P� <,��Z#�1����u�J/,��.4�"���.������j�c�K�Y�i��9W�Gb����U������:c�A�!�(匒�,�2���M?�%^��z��I�gm��K�N����p�L���']./�bRao��{����·�Ķ��V�׀��X�6�s�<�­�Q��:{�I�M�So�����+W:�/?�W�i��K3ꐬ��-���z���D��q��+4k~��`{=�k;{7A
�Ä'���s�}���m�����:V����s���H����׏[ֆ���/2�u�:�b��ǔ�.��7۹UC��-�s�N��� /�����	�շ��AW��ux�#?Mq�YղO�㸵ү⵴��U�I�
��X�\��U:	���e,M���+��q��w���V*��d"���a'��C�C��I���H�t͆�w#lv%J��*�!]�`{������&4���cj��c�Cz�{~�f���~[^��]��T��U�@��ȍ� }h^�p'd�ul�j�\%8f
��Z�[��Khbei[zpz�H�f$�	z	ecB˺��F!��=)64�G9���)����in���ڢ�td�����Iv��6�PmLQΓ��"as�m�bY�/.�)[@�1@\��%�����ʨ;<�0Z�*|�� }U�Ī��ɞ����jAA��c�!T�	�Pd�:?#�#�>�kNb�[J�Y Y�8wo��ݎ'x��8��ۇ@0����lw�������@��K����/$�`�J�yt�΋^��`�8⹝�	Ig;��	 YE��]��;��չkw���R]&q���Z��f|OPm��ݠڀ�l��WӃ���kՔw�ŧ]W�a �Ep��=v�l��a}^��+�ղG��0
.2L���"�>@59���K�����UQ�-���W�!+��Ҍ	n#�߳�<��m�}�g����4u���Pʺ`�Ai�j�ӭ�d9�jUX��u���ߑb8���*�W�˙nuG�b�T��.t%&���fd= &4#5��:ĤE_�=ĸ:ECsF�׫�Pi�������8#����mGbj	����i�^��Q!Z)��TLu��'�wj�ԝ1���{�B7*y����l�8]� &�$�u*�m����mrd�֭��1E���sP2AZ#%͌�&a�^�{U:�%��i+��<"D�>-uw��>���-/�8���H�Ԏl�2Xˆj䴧%������!N�Y�q˷/K�����Y|�>ѫ��c���:q���?�i���
JiR��\�<	n��I܍���q����tyN��W� ZQ9�E�-�_��[�!O�$9�R�Yz��B���ߘi�1�Ʃ@5?Ŏ2�Ϙ����gF�Qg?�U>��U���I����$� �y�~�fk+�tZ$������2�|�V�A��FE���a�AS�w�LJr�_8bV���$@�Ɍ������Ԩ�.�ft�ٴ����_���?�΅Kd���yæC��4�$�8���ʫ4�Zi&qLS^�6�h��J!��CG�Dib��_>g,�X@8Mu����~w����ޮ��$�aj��ﰊI8��I��Y��k��1��������*�S���%i�6|m9�����aє�}V�^	�[ڗ��IϹ�t����x�(�%7#u��h-G��X}]1Dqsv��qJh
��?���*1$�cu}�kܻ��ZB�4 �vgXդ��2�mE���i�G��9��2F�4b�_�9��M/�j�#m�jP�M�X��w$�ě!ur;��U#�R�] ���k��A�t"���G9���#�%q_��߾������C���1(�E�"��0F�R�GFe��Y>�f;�t�����g�&~��/��k��0d�M��I����}[c���K��?^+�� �x��E��܌k�*��\8$)�e5�����6�M%9ɉ��;k�Ɯ�Z�*^ϔK� \�"z0�x
"���r��R��ǛJ��Ԣ&�g�L�N�v��$�Ȝ��!�Qh���a��aCǔ���)I� �ө��"~k6�4��D���p����F�`�C2��)�����g�@�Fc�E�_���I?ԇ�0Q] ���0�f����F�{��r�)c�\#xQ�8�a�!�CȐ.�z�sH:A�`)�ȡ�n>/"D�.��g����+���o���*R9f�����Y�e6�aQ�AS�١�m���8��fg4���+N8��%鴩��� �����1X�Z�4�qZ��}ƀX��:%���۟�<R�-�Y����w�?��ܴ�Y��?���{�*�A�FJ���h�,���b�+ S�h��>A�>�D?��@z1�c[8L![�M�{�h���C�Z]���D_���
�a�ݕdz���!J䜂}TY� F�k��c�|��"�rP#�o�s�[8��_��o� /.ZMd�Q ����=�y~~'�X��
��p��/�x���(��Ɠ?:SV��.��6�����s Q�D�Ji\��r�]��A����u�ǪS�m��٘�t��*�P_n��;,�|7*�s���i���LK8R�V�2���p�n�M����WƘHϭ�=�f�n�� ����n�0r�"�ҭ���y=oj�O�!���j�R� �x7F�?�qr1���w��'�n[jG�*�.S����$�w�Ν73)?Rӗ!�M����x�=�����U�]��S#,���3�y��^�*��}=�j1nf����y?�6�xY��V�.3*.]���2#���2�G�б �W�����*;�Iu�!�CTٶL[����N�M����r��Cq��79��v�x��^�B��o-}T	��o�g�Z��C���u	�<R����6����q��������}jP���]@�f������Z�2��voy��^EYS뛤�5Pɇ���n=v�"	(t��&7�Ui���w|���)�%�i<8�m\<͇�L��r�S>W�+��숏x�SɄ.O�RE��hZ>:�wfu�К菛�Lo13�D��q�a@J��� N�,�-��[{���d�~�-���R�KL�nh�r��et�ez{#[OJ��F<4���-R|�^{��@ew�w:aqR"Aќ�n��2����0����v�(5_��V�Du�m �  ���jS�Yq�F���V,(��%2�ޡ@��,]w�=�m�O|6�f"P�Y	g�Y�%u�#�m%�v�f:�Y����ԞˣP?���u��2̋���\zk�)�������o�t������[>&�*w��r�C�fe;k��є����y��Wi��b)�_���ѥ��EkBܫ�Fq	yڮP�>гbէ��E��;��^��wi{��o%��5���c��C�;.ƭȹ�k�|$p�5=�P.���������t9*�����\ �p=���D?5j�P����~�#����D"����8&dr���J�chI���y�&S�?n7���V��^��ivuBf� zAB����v�;\h�U�+M['.?�bM����2�w$��K����|��G�����0{]�9�2��Ab��cg�_�o�_W��'�#�82���S�7��q?̺�M�!�{��=��ۊ��G��_�^3o��MrE��FN�d�
ܪ���|�[%Pl-&3��W��i�Z��kS��j �W<E��rZ�=�d/�InFx�&�1`s��R@i����>Z����<PJ��97�t+N-�Չ��������4#�_ �"gr8kU�\F��Y�N��$����$Dh��y�|���4G`;x���f�}&K�����X��JMm�� �3j3��X�>	�#m������1Ǩ�:�z�z����Suy�ը|�ܵA�F�#3�� ����>��!'�����F����|��&u�&�p���e���$�!�U��CWs�PR��0"�߬�s�:�%�8.�b7��o���R �7�,�w���eeLZ�O�ƩetR����ɧ����O���,���n�9��@�"-AX.���:,�s�AҠ�
���ǥ��L���Nӳa ���4EE����Z���� Ӕ(�ʲ�H���:�� �VZ/���#�Pyx	�>�x�����z[e�<#B0��.UH�rhȍ��,��P����e��R��N�i�0$@�<���s ����y&�e��	��cP�`4'�K<!R��]�\��)������ �!�i���v��@������(t�
�p��L�����2ã��.�B/�#��x,^�/�����F(��^��X��E�0�*2@����]6�Z��lz�:j�:�นn�@�%��%��Z��&�P�CZL�%>���� �'���t��	P�*DoG��H���<LL\+0Q����2X��W���>Ęk�{*ep��=w4�G�i�71�}�F���7\q��'Rs6W��췚7�ɫ�x�K`ŢP9��9�C
�0�?�z^nU׾�4;����v�C�����,���3:�1xٞ�}Y�r��<�2-����z�DB��)�r-�o��μpg&��CW�a�R&K����U�l9nlK��V�b���l����ڗ�uF4��#�[q,U^xhF���ro�|�Jd���;�<��yJ̨o������@)�<LQ�1��5W?�7�����CU�o~XN⹣1(��TWk����"�ik�QHs����C8���{}�]Y�0�b9�E�c6sNBt|�1.��Zy��N]��Qp&fl��}������.��q��ԫ6]���v�檈ݑr����odZ@l���+D�N�s^4S+��:���@S��9���|����U����<ʒ��2F�ܧ�����}���U�*�CϠ��;RǠ�Y�M�#6/1���ٜB���)#
��r�� &����$������E����g�!�#�'�����΢�ɷ$g��PQ��w�UQΨhs}��V#뼨�҅瞐�z˄
����C٬�5ń�5����`�>�Nׁs�.�ki�=���j����L�Ͻ�ew�J�z��T�M�͔�2�2ĉ`��kٮ����jw�M(�y]��I4S�UR�/K�9��`��|����l��:�PfIeb�~�t��*���ߵQ;�^Ҥ�_�t;�)�%�>������
hmBE�y��?~޻�]n�Do�\�UT��CTF�2>yD�����{.x��gw7� K���|�A$Y��Q�l����Q*( �$ ��A[1�H�U�U5?S�'�d鴌DMٛc��y�Zȇ=���6b�U����B�l�
��,��ب?_�����K��Y��k'��m!v�#ث'& ���K}vi����Ki	 m�0ZT�a%����"l}r|3��$�Aێ��f�H�W� U텢sƽ��[J^�x�a`��E%��9�|��p�M_����E��H{·"��D��ڵ�P�ub�tA4�@��ȣ��L��Pų[��3gv�</n�mT
��ܿ؈Fh�G�o4������l ����ֻ�z�X�0��wD��R��)��[��'�_?@�j�����t;��⤠��o<�0"��so�J�5v>��ͫ���=,�1ʠ(�X$)(��D$�	g��ǐ��Ɲ��ހݱ}}k��pqZ�G5]�!I?̒ߖ�GP^���9�ȍuw��VT,_6s!
 �y��"J�4O㎯yZ�">H�n���k�Z�
�)�7Շ�
Iť&�Ǣ�9*c�%rMD�\9i�bPC�w�<M|em��6�;��w<��ʺ}B���
�tsr�Ƅ�����/���Ҽ���ÖK��W]�5���o��)�'�5����Mڵ_��Nj�Jt�Pb1�y.�̽�������p�8T�=�{��iU	V~kB�$A7;vWS��{3[&���޵]���[�4�[�)���(|6E>�ի�����K�$���V�A�	E�#�ǂ�.�����":&�_�'%�]6-[#����d�?~Ѡf|��&���d.b�M�$~#1�G���ذO,�O����$%�`�(S�̣Zc����3�c�22N��J����6B?oC��Uzi3,{�'���	ݱ\cg��/9z� w�W"J�E;~#o��%\������$W6�78ؽ��l
��Ɲۇ#*�X�l���3�W`�i�4��j58W��ͶȄ�������Į&��9�^���P�5e-�B�7
�E���}��XM��`z\1����e̤���������B�!������]Ư�T)s�t�'$��wS��ˁ�M���I	�cxm�+�H�oy}��D5���8�oi��h^��γ�S�BU����P��#i�������3�k�Ɂ�+u��o�X��֎����D�o��� Q���ځ�D��UǸ׍k*��(\`F�k�vFv�OB���A�U�͌���G���ӖyÏ��g�~gs���-�8b� [�F�63��t �ı�����_�����,Q0\(u�7�c�+`S�G�Y�l}"�4�ҫ8�~f�86���\-_�kYNІ$��m	*�n54.J�L�2
I'DH��hI�,��XA��򡒾�Z7�S�&:ø�}�Y�Q����B���s�f{b�b^t���[��$�q��Ӕ��F�t[�=�Ѕ@�����So��s۟1�l�~��C����'=@���8��]���fG�\ǌ�o�iY\Ru�����n�ˡK/���ٗv@H`��Br*?��1޺fo�ς��;p8�����{�����ګ����-9��ȓ��9������8��_��%jC-�E%�:!G��au5��8y+��]!���,��I�X�d�4NU�;>�au��*m�H���r΀h��.�<%�U��C1,��;������������A�|����22��_]�����c{��^X�hخ���5S4�Ѥ�O�Lb��������p�i��Y���Z=��[���\ܘ�,%�yE�Z�c��Ҫ����J�=1^l)b�Y~����W[��b�{B��R�0��üz������I��U�Q�|iۈ?�1;�lI�>��ů�M=f�{I/x��i:�..����;�3�ZSkM�@��C�c��A�� uq��R�` �Li�P8���6���t8���ĳZ E�o}<A]�.��j�Ů�-�M�$ �`��-,A�^�EƓB��b�$�<fX4+E>�eϱ"e]�$Z�֊wQ���E�l�`~J{���w�NO���|��!�������4k|c�	��w*���	B�� W��S�Ҋ���!��Z�8@�R9�{�<��s�0\�!�*�7>&�U���	W*�^�>L΍T��O])��^��x+���w� Vǳ^KŔ�Q�Hh��U��y�r��"s#H�h����<V�߇@��6��/�yo1��=G���2#�[�j�M��+Ή�r!?EQsY K�;�D�bk\�tH��P��5M��;P`,e?�}g��P�L��V��t<�������� Ev�=̥Z��;C6�D���^���#���<i_���C���WD ^\�s(Nz�s�$����Z��]�2�@xdD�EO�1C����nEW��lt�GVD`e}j��s��w9Q)6\}�5^�m�'�gk���7�L儴*)��hoI��z�uj
��o���<�����6B8x�N�m���t�b-��$a���jud�����nuR�
��:o<���R�*���E4R��vȩJ([R�	������C�(����٬~(#��SE����U'�W�	�뮀��k���G���jMո��z�$�A�r��B�Qe���V7�'kn�P'��O�)�9~��!F�+����9:�@�7�"��"�l҉j�y�l��DK��qHT�-�hBY,_����!�����~�&������~ΐ��|�<�*�Y�K7�`�C?_N���K�e�^���i�6���O�f_�y�J��n���#�Ǖ�,K��5J<b"9��#qگђh�޼֟jӮ�hgᴵ�[���넥���<�E�A�����F�B�D���^k>Ċ�+����KX��:�D���ׁ�iL����ky��������Q^X*m�U:�����	~��메��'��ٸ��lA-�� J�\�4:m�R�&uFb�s	K�mNf���
�`��n�Y����R��e&c�~���Ȅ<���4�G�׽�.���Qd#S���hq��a쾌��,�<@����k�fɬ����$޳1?���t&4n��ݞ<�-�T���_%y� �Z� �t-ym�k���o{>D �f��,&���̋���I��.{����×dRӿA���@O��w�W0W	�?W�Ö^���EĪ�����Kk� �,഍�W�M�n���n��Q���*K�����i�D�~�.4�>�X�^��.J���j#��SDL^o �ߺǱ�=�~�=[jU Ѵ��$/[�fz|qZ�Qv:M:�)�cRE��s�<���:�
�&<���Iͺ_�}��z��3Y���`:��,�v�n����������s������J�k%8[�IMO�$A��a�q�;p���x;���2o������Ԣ�B"&(�Zn��-�",���O�� �O�y�$�0���O;���-=�5�[B�z�P��a1uf���&�J+��Ap-�=�;����!+I4�y&U(���b2XZA��2����1��B֕�@�<c�]�XU���cV��g����(���;��^6{):ͮu����t�h#I(���سz�;^�W���.�W��h��+ų����^	��暻G~����{�F��#E�����f)X*t��·̈́%����A�[���P�-uRԶ5�o��ft輢�𒎓��f�JyE��YW��cH><M�3�99H:� �~[����^�mJ���C��������
�Ϡ6-4�5u��,�W�敲���4���$9.����vա�).�W��[���j@�U�֌[�O�������R�=�R�=a��P�b��{��g��O�V�{��^\3]�3� O�V�A�O�v
�WT8��골����1�z4��K��j���QYri����I7������G0���2���m,ʯ��� dq'gz���G*�a����
;�v�h���!�e _c����^�j�׌}���0���^!��7ow�J���XFm���veP#�]�z��1�r�J�5l� ���y,����������ˎ#{�єٯ����)Rd�X1d�Ƚ����k4H��F0�h�l�et�C���F�� ��@��d[�^6�ߟ�9�ﳖ���cm��V&a�D)v��A[��j��j5f1rp�>���>�[��q�=��)�Y�FX2�S��7������ȼJ.g�Hj�pLi�������8�Ӥ��E͏����m=/�k�����)���ڼ>������MtK5��1һ5���\m�}%?ݗ/�JBS��T�W��P�9֔�/�{�D���qD�JU���¿��Y�bQ�~g%r#���Ob�v&r.��$=n�;��*��*/"f����ɰ�_@ԁZ�9�_k����a�QG͏g���b8�T������'�Q+YHbb
�>��/4����XC�^6{,��V[.Z�V�CBmK0�n�������Ǳr<�\�-��߁A�������yO<�ӛP����Ƞ�6�z��|}�"
_j�O��'�sONE�5fJb.h�5^���}]Lz�빓��T�b�HVk��ٲ��L@G����r �1���W�E.uȻ��i��{�cL�:��:Gb�Wr��S'|&s��X����yI5[�3o�d���S6�ַ6�wa_[�'.O�p�֬�i���ﻘ.��u��i�Jq��>4i\2$��;�)��'iիBԪHc	ɿ�����s�~�"�D2���a�L_L�G�M���_P�U���p=_�²��z�sYCb=hj'#+EnI�h�⦤�YkC=L����τ���5Z�HU�%,�K�j�ٕ�"��Yd	��3�8�M'��mN�VC������G�ptdm�;��cfj]�s��I���T��A;"Ʃ��?v��z y!�����CFȞ`����/}���Ɓ���eJ�$oM՚0����l}���a�!� ��*�䵸��Y�L�"*"(7��!r[ȡ>��w�\�~{����+;��Z���%i�|`��3$�ʖܚu�0!���X�]���Qz�-�~�Q/�Ҏ�*�D*ߡ�Aj�&��gC9�ԥ���ˠ��.�K��/��{ E[X};��b�f��N��!� Y@f�,��Ӎ��୤!(��b<v4����*v\�
/����ca
\�������f������$�R�M�aH�����Lϕ}��2�+b�(��>���R��hѯ�z����w.{���؂[;�7��@�n��Z�?�2�Sw�Wz\B��щ��Ex��ɟ�d��9e�͊�r�%١��k(kkz�C���/8�߼=s�:+�/C�'�c]?��#�ޛS��p�Vׂ�b^f�J�35G�ĨFL��2�E��p���$5��d��N�׍���d:�EF <���;�9������DM����>m\�Q$�t#˔*�ݫZ����b��'N.QUF����dJ�1���4E���̢�qd���뤁��V�qF.�j1k�ZE���Y�8��LJ@�X>�e�2���3<{ﰘ���S�E��<-��B���6�N�����֠L���$	�~�1R7���@�ǈ��:��|��ڻ�cc\d�B�5}=g���'et��j��Vq�m!�b�Dl�H�qd�S�k4��%��=�t�H��\e��a2I�(�y����\o���q̆6iB�xk$[����WW	�'��>��������*S��I��3C��1�E9���|��g_e�/�*s�:ҶN v�ٷw�o�����Xmw��0�3���rF��͵Sˤ�xu���1��AHJl���sA];=�Y1VD�R`4�V6Yu1,�.�s�7���KL�Cޱ�t4r��h�T���݅o�������,�x�$�B"���G��S�WB��d��]�1�����Z9����p��-�����55�ڶ����^�J�$�Z�V�.�mx$�R�kM'��wC��`��Xc�d�H�b(���±c�J�a�a<PP�F�/]� $b�����1Q�ǫ�R�߶�c�Jb&�x�_�`� �`��Ňr<��k~KD�$�j��ԯ��9&��~�ċ��$�H�.�1��M�����Ue6��^S��d�8>`�\�U��D�;XOS�(����2\�mҧ��C�$E��R�toU䃼iU;#�'q�	���¸A���s�e�iq8�uUVH��'d�Fi��{=8	>}M���1�=pH惀Xx�oQ������O��I��y�c�_.mz������s��Q��~�v�����ƖK
�Q��x���x3i�
QF#������r��=�L/֦�,.:"
�=���6�?(�JS8<�}�"�$�>��O��ۄK�w��LT[H��[�Dqn���T��2%�c�9�n����"Ѕ�1@ʽ'��Q��#[���0E��a@���bXq�8�9ωM�t���׌�y�C�L��>���A�R�K�1�W��l#pG�:CPh�9{tbt����6�U�����o��ȧ���C<C�pN�ic���0}��>�H�3Ap1����;�bk��xw����X�.Gp�c�x�]��h��*�ԩ���$�ώ+�Ji�^O�$����:r���mY�5��(=z�쀹��nȟ�ؓy����̤������2nv�6G�q>��b9u��3�9�`p5�	��~�\�6��� ��2�W�������Ԉt0�#��Ј�q��	N���$�6\�k���>vK{��t��m���`1��m/�]X�r�6�C�������(=,5Vd|�w��X(���}|����F'���X�P(������n[��p��X'�>����5�ye�xaeɟtv
(�'�:���Q�&L��q4&J�L��u��xP��x�>��]�dױ��w��I���Ȥ���70��Z�w���̚Co!�������+|:���t��}+�۩�7�[UH�&�	s���<�n^
4wk�怞�gE~,��J�qN��9�IP��9*�֐����z7�QGMpTAm�#�2R�4)�k��6p�~~rӽA*ge���3]���
ї�]z���HRr�Lx�N��ΎPB^��XGʕ��F��I;�6�逧W:x���1c~u.��Pa~��"�Qw���/�3�|�A�R]�@P~^�y�|�����Z	�~ʙ��Ǉl�������-���0�6"��J�unR�<�h��? �s)�"j������'�;��>�K' r���H����L��=��$}Ц��p�,�A�W��}[�0�'�ƯF��Oߊ&���XGɊ.� ?�}@���y��=1�2�1��O7mY��D���OBpD?���'nW�?����׆"c����?�[�DS-��q���o=�}�އ��o 폩�RG���{�@�Z�~�t���k��e;��uDR��������/3pK��G=��oڔ���e��^�+�1�A��@�V���@4W�p,�K�Vq�^1�5&yJ5��Ө�Wu s�"ҘO��O�۸Զl�������e1@�J.M��\=�6������;"��η!�uD�w ,�����D2�֨|D�>�F8� ��&&t�n��#6Y݂��Wk����"]ѩ�-f8��9I���j舢^%055����(c�^g� �Ny�q������	{�D���K"�ǎ�eˀ���m��"|���QWI�c�tJd�Gz\��E�Ț�p�M��R�9������<1˻a,�-�l����{�_43$���X:�^վr^A;���'���p�{�v�pH@�{�[�yS�)4�������T��Z�
����}J��$���M,����Ėە�1�Mk����L�[:�qϥ'�"�8m�{cf	��Tc�߉����GJ��.��3��]v��h~�@٘���ۯ�rֶ?}�_����UˍY�,kR��V��n��i�^	�Q��Eo*�?8�G<n'�j'��$Ԍf��I�̴�����K}����V;�#���&G�x���x�|�3s	"�O�m�d��^`����'60>W��������@oi͡�J��rH[&�g�� ��I�}7�}��)7a��6Ԑ�K3����א*⒡AY)a0�u-**r<K(f�����w���L�C3��ȹ<�NS���$/����(ڣg�&gJ��u"��:��r���9Op�WQ?j{%v�ۆ�s�j2vԨ�%�� ��X�9�n����Pn'�Qj���ox@�F!U��g����K��0һ
��(o;/����S��D�����"���hj��.p�d�ҋi��gx$2
`�`��8#t&*�M]�X�+��N�������N�~�}?m:nX�w���ʉlX�;1�Ͷb\�fuH4���Ɔ�Y�T
g�s�|=�ES�RbEs �^��m�i�4O���e+�·=��[b�./�� �)�8�`����I�mϟ� �EmOm�zs�RK��M�2����}4�MĬD��}�V�o�:����;�í�8�b/OW���`�"!q�#�<����̳Z_MY,��Dp�KX�x�JV;��df	(�e�0�X$�9-�������1\0 �rҪ^�n�I�|�Zs�����q����QB�Vs��8�W�T
$���h'���"PS��T6���|�0[�z��C�`�fD�ץ)�i�#�ًp<���3�6����=rgZP����Y0��3��_�E�{%1TW�xU�z:�K��nh�ö�J$��c��l�"��Uh``�v�T����k���u�<���?��D����I����uI���v,L�j`�b�#@������������Ɂ�5��ХR��� ���[H��W�=��O�%�X�;����
<�>X�o��D1z�*��{>�Ə8T��'M��U2��e�x10.�w��1��x
�#whk�=k�	����+��U�vA�de�>�����O��xh����wH ��y?�k�����]4)�,�c��V�:�2�XA���4�v�]:ʺ�����	Fe�c׫+�����E���ZO�|���q �nT�T�>�⪮�P��T����!�s=$(�������C�j�h��@���&����u(���:�D#a>1Q6ݠ8X^�#�GL�S.s)P�;�B�E���t�Z�ej����	lkK�J1g{����&��!'�)t\�zdE�b�-6��9��KW)ޚ�4�E�o+j���ji����$%�<��5��'g"sE��.H1 Jl��Vb�f6�*M)s^}<{^��P{A[�q4.�N�
B\N�I�,x�4���G����3���������/�]�>U�-�ǩ+��6�C� ��~c@�m�m���m`�3�5)	�,O���R�t�w`ՁߋOG�Ak�`h�u���-~�l�_2��g�k���v����)Ȋ*;m��sT�_�k��W��c$�/3�"�(ܝ���~Ͻ���l%*����0�f��y�I�3A+�\�Xa?�QO�ܓ��L(���O6�kw(����b?���&����W`��C��@A���VS���<�m�h��6} GrS^�H4��,�~(D��]c�#]��[�Q��*BHy��f��:���p�y� "�Q���C�L�i{�z��i�+��ƥjo�K�|�ۈ���t�������G�t�>����V�녻����,��X���Gν�:�r[�r����̴��������˼������L(�gs��WNB���%2����>����
�����֙$:;ZAQ��KP�電�)�<��:�Ӣ^Ƹ�� �H�������Ο�+�D,ה+:�I����nvr��o5~��cm���pU(ˋ=������Fd�M� 'ekx�=�v����P���u�a�����1�L����b6��E�;��/4�zx'�e�m���� ��R��{�n|Ǌ�u�V_- 
Dꭡ��9��:]bk���;$�˺I���uWz(q�)�ٯ�-��裖8����x�zG��Ҿc�Ѐ�?�Ji*�l��R	A�O7o鎹���_T�IjqI��'����v&Ӂ����p���0}x��a� ј�Pw^<���
��WH�BnUs���J8��*����jy~BF�vB��dLXK��d(�ˢ)\�02�U�X� ���o��a��N��$���1-,p���tfW.Z����dB#y����f+�Jt�����d�a��}s}NeȄ��V
}��IlqZ�qY"ސM�]�`/fF.�B�=�;u��Q2p,B�'�X���?�I��Zw��]�*KY�p����$�6�D��(l��eh��3r�~�=� E�4^ �G�������Cɦ�c�(�t1��"Μٱ�	"�Y���nP�M�.k\-6v�Bs�w��dz/Z��W�FN��SrmN���S�����؃%g�$�%V,.�����g����ℸ���%Gx=�^�u��w_�fi��,��K����vCS|���Vʷ�BsY�]�R�:hѹ�5UF
��4�&f�6;b���nV��?Y�lOY:�j8���$���Q��j=���#]�Vx3ٰip�%�����9)����7P�3�ږ}MX!������B�v�,h�iH[B�ޫ`�����=�wY�+�瞄3_��M�O��Gjjd�������@�9�c�us�[c{P��&ƭ���(踍5^:5A���m��	3���r���D�zn�=��4�Us��(19j\lwd!�\���aF%��X��;%�,ed��Z	,��	����P'�
�5�;)�8ls�SH\��6��Pu�!|a,�2���.m��F׭��mo����67���X�a��Z9�%�y���m�Fy(�;���{�w#�JB7a�c��h_�ߙ9�=D�/2~�,���pG��Q���c��}�F<�ûv�Ȝw�4�\V��CRZ8�ț~r�g�{_��d?`VQ1E�η��#������)�0mth�,�s�./�Z^�;n�g,`u���R�\����n
�(��g0�ש9�T�{WaDS	ֻ�bА��V��,�*����ﻓ�����}���������M�
��U�xއC*�D�O�$���	��3��܉g`�tH���H˱TP�]G���Ӏl�Ȧ�Z�u���S����ЎM��ݑC}��)'}ӫML�ĺ[�4b�eE���{ҵ��!Q��+)����:��M��x��'T�� �Y���2`����pF׃��mxV�q#�xrRe�xyXi�M�Ю	�W`,
 0���֏[l0&uRVc;���@X����v�KZ5TPr:�gqw���?S��,�g_�A�+3�R���z2~�4��JM�L���-3�hE��G����a��0-B��Kr�n���2C�Xpo6�E���(�_�pr%�J��t�((s�xn{�%z!��9�@�y^��K�8Q/+���>��g��E>���Kj�A���QLm�|k���1�o�w����Gs1���@0�������ĎRO��t��,�g���D��T��ԤX�=�*�b=��tO�ɒ�dĤ5�D=�����lȃ �z߬@���fVR���w�Mv=S��[�9��G%���$<0�8פ�\�E"���V=&vG��8�WHZZ��Y�r�S�ڶ��};�Ǉ�S>{�ު�p<�4���0�R�/|��+Hly>���;��#@��Ĩ�?��y4}Q�}�`�������s����B�B�NىT�Y\8SKSn���3�"6���������]��J&��ʫ�p;L�k�Z���W!�y��WU����Z���#%M;�TKQgg���m32*e���ɹ�=WaԽ�y[@I*��q#�r�X�����	g1~��.����o��Ë�U"bn�"��H��!�o���ފ��2�/OZ���r���;Z�[x�O�����R��d�o�i��a���Jn]�.!����Ws	ļ��`��eI��e�哛�a�/u��x�)�5�^/S��yQ��|f�$`sb�8A) kzT��$�_` �r�G)	�ꊏ��o�g�e�QYtr`{�xM-�V(�^�{�zX��K	ۅ(APK�DD�3 �%����8ÿ��+oTO(�7g2����9��c���C0�]�SnI�(�3�ZMM�.�LW�ǈЀw� �j[�mY�����]Ҩ��P.�)&���Y�:*{k#̼;nn�=0���"-���v�v+�>����塗6�z=U��3T��i8���>�ö�a�p �(��;J�zhch�J^x#��/��1@^T|E�}�j�R�{���!_z�ؠ�r���,�y"���į+�6��YT&ݬU��ų�j�p�1'<>7���\̌E�
�)��93��l~��U��m2w3�=���2H*Ӣ�-1=���	T�7|��߯­�h(Kޤ�>����ό]G�V����"M�xo�[�X�g��������:@p��F��4��ڃl�T[��}3��
?�ٰO�nc��U�Cޜ����_ҳ��HM��e����{c"I=�S��� �q��]���ɭ�{Ε=�2�,��5��lR�ʣÁ��n�}vZ�%�E9a&���`t��9����fz��/�P*5�R�q&�?3.�+۾n$&+���j)-����9�������d��� T_.��=D;�~Zټ�
��|ǽ��;e;��R�@�#�Hg|�KS��Y�������C������Q�*AF��L�V�F��'״��0�0��AD�O!L(V��J����hr�l<�r;��u1go�݇�{�FA�A ��N�3�������f0Y)\Ƕi;h�-)����2�y=�φi���?�AD�� Ì�'M	��ZPrH=<�eZ=�at<`��[��C;�N:��ZY�-�#E�<��LP�60��$���{������wr3����C;������Üx�~r���a���O�9:���?�Uq�g�ꗍ�2'6���*��\�?���OR�0�����0uŘ^ԋ��O������ǳ�U ����L{��I��Q� �b�#�������B)�pVl���4�ls�.eF;�"�R,��b�߶���▔��һf��qwmQ P��VvD����TR�>>(��-�\��G6P���tꆕ啪���һx�N����}H�(@%�FU묆����ȧ)��d�y
;��Ȝ�zb>�����9��=�W�wt�¡���8M�Ŵ�K���@�0%։b0���~�A.@Yԝ���T��)�j������;B�.��f��+����3�VEK`��r���?�R����Ӗc@�@WV
�^jA�ܹp@��*��z�j*"�@;�O����+q`"1�y��I��أ#�]���4�4��� rP����P\��/lO i��<�������h!� �u<5�9��A�[���N7��ì�nT��٣��q�m>kG�!-o�>?&ᆗ������M������J(a��Q�$�	<�A��6՟�ڬ���q�*I:��lDH��FX��-�⤽�ĺ1�=JRG�DӛrĢ.�U�5��֬[}��Z!�U�K%����깔����kU��Y�T��+iqh䪟a*�5됽�qYm��OZ'�aT"@{��j���z�����m~�٫ײW3��Xl, �Iy������d` ����
"���\dՕ�N�ɧ�e��ur�ע��º��K���@��b')Y���k��V?a�so�*L�����0r�mY���V��.��G�C�cu
%P97�� ��'�����_�;�~D��Q�6�x�Ƶ���B���78s����x�k�`�`�%q���������������+چY�G�m�z�΀���o��H�w۩�q�A�"�y-V�'i;C��ꨂ�i�c�u���f"?Į����\���_��4գioIg��
M?+^X�N��8�Ƽ��@��K�9<�\sW4�����h.��uqa�>:�=]��F�f]�� [�C��̽&���(����;ȩ�e6���������p�pR�Qc��Z�C3�\wʤ��+���VO�A�<o��X�3��z!S��Ob������πW��r��Wȭ|}&��"e�/Np���w��né�4x��a�]Z̪b5�%�$@�xt��;^���s˩�1�HB���_(�z�rs�d�X&��$K��nF�_w��A��U`e�T�w�@�P���<��#�a����b�ˉ����S�|�L6�$��{@�g"�U uL`kf�}�P#���<�D�[�V�X���V
ܠ	���~�����o��p0P�~7��P�� L?Kyr0*�:%��Sq6ꠝ�÷@:�r�X:�N���
�P.��!<��J,a� ��V�{Pgg�'�=�N�)Dg�ª��ޏI��m� 2We�g)C���V�A�%)"_Ӭa�_z���;��QA�0�2��?���L8k��f,��P'67��H�BM���6ew>���Z�A�\nwq`���ʐ4�,��l1�Uɤ��Q�\6vg*�EC<30�T��!�	!�0��ꌼSv���*��eۊн�,�6��T��ɀ�t �E)�í�{�rL�J��{��!�j^�ۻ��
̾A�F���hL��jj
���a'�a���xIF�Nb�R����@��ҎP|W<�'�Q����Wk2չn��/�:�2] [��V�2� In1�� d�HY��ts��b�e�H��Jt;3m�qI�Z2:}�����/����qB�£x����-�4�Nfn�
Ɖ}�~���ߙ����ޤ�Cz�yH�̅�Ul/'�u����c)U�����L�aQ�-�RG�H�V5���_`Uؤ�6��@�JH}^��ܪq����1��_�\�n���y����w���3�7o3=�|P, ⥌l�8�խ�����&������
��S�W���l�$W��Y�!��'g�*��@�	JN�0�Y��c��%Y�C��E�� 'vTu��@^��7��q��� �h�����7�R�)��@� ��3~�Z����rww}.]�I��m��q��F���@P��_�����U��*�n��7����Y����!��& �qa�!�A�����Sۋ���j�Wٳ��&$� �/�S7g�S�xTa&!v�������ѳ��k�DJ	\�ƒ��B�x`%��*
O��[h���x;A������4G,�5�ւ򉭇Rߺ��w�s�~,mmf�\����|$�i�����u��(�����^b�5�y䶹��ҥ�0��(TK`�X	.�K�V۲m��&�H >���)G�:��6X+�����
��\E�i�"a0�2_���֓��[U{��'���r:XU�m{V!ݿ���POR�6mÓ��{9q!v�;�Pu{e��t-��L}�Jm�l��{
Y0���`7&f�
cY	P-n�|�gZ�4o��P_��������:�m4�䒙�*%D������4�=ˡ�o������h5�l*wG�/e�Lȿ؝�Ԍ�z{}��n�{��*$�}�e�t�J�يDbs���[#���O�e�:��_^�7�[��'f�"�|�9XQ��jz�/Y���0�͢l�y:�3&��s�1�S��,c�h�G�)�$�|zܖ�7��e�hOo���������k>m��x8�-�F\ᡑ��b��V}<	殨������
-��ꪤg�.<_��y��V��)���VS�=.�@�!�9�0�aٻT��a9=i����д
��L�w��]\А��mZ�.m��v�������
�]�a�Xf�'�q{�p�²�����q������M����lɛ.$]  Om@؇>�+k��h�G��(��H�|�w�?T@�A��'��'o�1|����C�Y�T_]��0�(�̃���4�Y	�E���/�������p����)x�T�@f(�5Y��O��� ����γ�8)B�m槎�6��e�Rc �:���e��������ꂥ7�;���R�&�kP���l��Φ�c��#G�wYu0�u+b?�ĄbE�]cE�,��P���0R�s])��p�dR�@�>��`�4�[˛��E��	�j���ڇn��S�`XrlJ7��#ر�v$�;���(�����R�0�X��/nZ���
�����9�NW#�j��.7�0m,q�)�dg�$:/�>?\����^�yL��t���5�z�g7宭
G4yw�&�sՈ�g߅A��5I��Q�$2<�J1�r\���xD�S!�����Op��@L�ϔ��1n��-�0�^���t@Y�!^@��b����a�k��G;vZ�PF�%������	.�٭�,z"�Z�n����v|���TD?�FyD&�T������:V���-���j\O� ��������.9�a�cPDF���gpBDWA�Y��6���ϙs����d�,�Gr�=j�VRx���1Y)��|s����U�Yt��Yފ��Z�%�}D+\Tn�H:�V����&OX����5ַ�H��i������#�v����.�WģMVB�i�L��0ñ �RX�*]��*���C9no���a;(�-��ēby�>g��Ƶ� �82Q���x����{��_ 3�.s�ޮ4m��G�N��B�f�wa�$����U����s��lk�O��|���g�-à& �?�-[�v�qӋf/
쵊10�1\���dZ�;���Uv�-V��0�z�X25~h��FΞ��A�������1���+�!�����o�	����	V�)��n�J�Kz���:�|��s�����=�!b��z�-�NǴ����pI�zOy�Řa� w�e=E9s?�sSjaa/c�tz�]��}}c��H���xLO������ׄ���A��u��_u�wv�D�>�M�O��-U��x�p�)�{GP%}��Q�	�|02�,�?i�fa�b� �R{����%{�}���<4�Z��c���Ry0�G�F�g���f���߷t�G��g�� $:I�Hխ��o�/l�R9�G��9y��%jA����g���A���� ��F�5��5ʮF�n��9N��A��C�c8�a�8���G5t�v�P���'�-4�/���i?w�gͭ�g�m�� p��7�Hh42�,��ܠ�=�zOi�5IZ���v���֓)�K��c6�Y��w/�����+�cMu)�x!�)����X��܈^ '�($GnU+�s�Z.���q��Z��&v���21���oFj���F�Y�z[�W��|�f�]*�v�I� �p%��)���@,7����|�X��Q7Q|
HC&C�1̎�0�{�f�yսm��82��m��r2'!@L���ܱ-�!�^����(y��+�kk}|d`���|�i�%bU�lCC��C4�$kRq���ZtD�g�@����[��n���,Ɲ��^�tn�����T��#� �D�O8�It������X�����2&�z��+����X#�"7����`�;Čk���Y���}��XL�2��μ�Ҩc�b�|F��l���eۑ�����,g��| ��𣮳�6SO��Gb��$��b!1�J��uVLԿIȡ�֣k"�N]��Z|�Q�yjs#
�.��3�N7�Ј�_��n�2p+,�4>��G(���N����G�{*�`�.��=[j����a&�Ш�BV�v�%�fڦ��h(�vxOT���,	~���^�n���X�-@���������~C$�n?��?'<,�4��8ɣ�޷8&�)��EzX�!�"��yF_���N.�����SS�\K�G�c�9N��vΠ�?�����M����Y
K"����Y{�4�~ʧ����0����a�^��$��T*Y���)Fd2�y�]�p���?�Ϊ�</��V�H�~T���FT�����4��]'L�*4z�O��~e��F� P�Zz��-D�f1Nօt�L#��	��2�{�e�4��`J$�����$zL�u����g�F���O-��0@Zb�Nށ����	�9܅R�@l����&i�LF��R�����y����/�>$w�MO<]sv�.�������nR�Eo�Ө�0ö��B�����u߃@����}��҈\���YϚ̮��IW�I�UV��LZ"P`���m�$/���*(�l���������{KJE�Z�{#-�R$ɪg	�w�#��F��$ۃ��s#�x#����Mf
��۪/.�a����~S4��M�'}(7#}�gŒa��-�Nt^��K(\Rz�]�t�Qr*Y����_6��O����=�e(���V�K(9щ�3�h=�갼��j�]@�_�=Qpd�b�|7�^ @8ш�ZaۿF�����De�i!u�Q�9]>�<XDK㽐��qH w��}-U�֑������C��B;��.�3����݇z���+z�9�hW���r��ǟ��"gEa�2�(t�Y�ߒ��C̒��0I�$��&�p���~A\��?a;)%�P�5�x��~��昧�(XuG�7ZftbB�&�#`$9'F�cC��2�������$�G�f��si�Z��4�mJQz�P�{�+�{E��t�*�T�}=�lO_��G,
�����������GɡE*iUV�/_���o.[�%���}��IDU���)1���oP6�8Am�F���n�tz��v���^QY��f��ԍ� �v+��ȍR5����� k�����r�r4��Z��"�b ��3j���UU[��9t� ��F'E���:fv(/q�����L��irY��?�HW튆��j;W��Fɕ���6�:��{EB��ù�� �tjU�ef_b;�ڙ�߂�������j��8<��ϑ)�R�����z0�"������7��M�f�:���L��(lKtY@a�����=n�{x UMʓ�K�B����t�3��Ɛ/�g!�egDd@�kӖH:����d-�WI*?8�Q��~���Ak����;�1Z��ZǞ���ډ��ǟ��J�w�ǆ��M3�=��]���7���J<1&T��S��S,v�O����-�h�E��{U��|�*��{ya|��p�G�6=�򘸀����[/���:p��.�5�^>�v�P�J>=n_�õǷ(�F�n�CX�}?/;�~��܍��׌�]�9�(��γu�>+s0��%ۦ��p�����f�rJ�#V�l�;�7�`E#E�y�DR�>�W�٤�)ɇx
��g��J�\�w�
��-k�i}������f��C��[��j(���<��6�!\���'���2�P�u����qsf�w� Z�Ip��J�Q]WMVU�z�xmp'XÙ�h#7S����)Ӂ]�c��F).�:`�2#i�I��Eq�H�g������\�����`��>{����W��+��H��`��1���q�G����1�{��Ǉ�e�KJ�j0�L�����&��������B�X����ek���/�`�&O��Dv�(Y<T
/�dpD�*�TҞAO ?<p\�q�WK~�Fυ�?#	�-z�tYq���룾g��hyg�Y�
D�� &F��Y��خ*{g�*����L���ep��"5B��%zl�ĈZ1�^gJ�)�W��d�.Ɛ�RGȃ��ى�Tsq�T��!E{���Fң�v:��sX����eF��#��}|��w=���|��UL1_����`բ�5x0B�o%A1��!s��ܴB�>��Ee�U94Z��Q��3XD�ܶ瞁e�S�0@ny��e�5�0�R�r������N��-'	OWg�^�=Q�4J��G�n��S��xz�5�l��9�#<mi�f� �����:�[[D��E���5��# /�N&��7Y�T2���;���G�)3b,���PX����!фz�93�.��	ye*�/8�	�TWޘa�r+,��$������܋/�ug�B�9C�3##�T$=?t:��+Q��S�y�;�,݁ر�5�L�۞��5�)�r<��;�[��$�� 8��3�c�����Qk��ƍ����b���E�{Ѿ.5�h����J�I���^����=ۘ5U9rT�>&#��Ü����bN�F)|��a\��慙bМ۪V"�j�k����hAƄ�p@Z��J7lj�-*��h1̰�9CKO��pe�&�:kS�#�� o]��,omR]�/��0�C*J�Ꙙ��|��4��Rpo[tO�'�ZxΗi-�=n�Ję��o�P���Vd��l�ʟ�3��!g(�)�E_Ü�4i���v{��?��Gb0O',sZiz���Lq���
G�z��q8����<b�T�-��xZ�b5F�����y�θ�Cw'�4pB�ܼ<��: :�ZzN$���,H/�h���@��S�{������ ��gҶMe�"/�CW�@iHJ,AK�����7��!�̨�N�8���E�iw4�s�Ms��h�C��#��,L���5Li�d���a�3���?�:j`*���?���o^�es`�=s�*HD'�\�1Ő��6�����h���㸟+S���YFq3xs��$Y�'z��e��,oQ��v�Ձ�bXU�j���cQ����z��'Og��±K�xk��Ӆ@�׶]/���޻;z�"߂�ˉc�LY3u#�7᪖����
ʾn�.�U>qe���b���(;:��&�?s����J��S���V��hF^7sZI��oH�*x F`Mk��<�Y�j��]�IHƅ��Ŋm����� 1�^�5����A��R�g ����t,�{���g���W}� �ћ��R�2��Qb��������4OK�kHD�b��mj�V���S���Ud�!]�� ������[�̻g��s����:�gF��ΐ�#eb�˲2O�܂�v޼��5���p��>��C���6%^�l����$��C������n�؈+�E_��Pˋӛ��a����#�6��v��Q��´b>�2���V�uex@�YƸ�:?��m*��<N�G���:���;y����6�Yjs�q|O��:ժl��quu�Jr�`{��{9��o`Ω��W:�In���hf
�t�������N�qظ����)�1돂P X�>0B��M݋���lb|6㭓��z޶���n�ى�i��=�������ln^X�tV4V����au!.�x��eD�V8���C��m徉Ίr�&�ztۑ��l�&cW�ª��#w���,р!k1
�b�����*4�s�>�5��I:7���7�'�a���=��?��b�u�9���=E߽0e�n4��T�#�S�U�v����l� ��ˇ�>�ٴ�� r��7�g[R�q�E�j8�S�yv�,���5�I �p��I�r]C�1�| P�� �'�G`Ml�צ��$���~0N�����Ն�Y�gf��n��&89�gE�ַ�f�&-����[��l�8P�zi���"��|7��@S�ĽA���^M�5���6>�|��xuWܗ

J�1��ʇ)��nJ��/&DX->i�~3�'�R�BA������n����]2��3����7�d����_��[B��d����k8|l�88�X\�Nߟ%�����_@���'���l�����۪��Fn��YcD�'t��qie�P��B�����W�-פ��d�ٛ���T{�Y�s=j%��y]o3#�.��>S����Xk�)&8�RR �`9VFX����+�f�t+��P�I�dcB+*�M*�O���'�X�Л�\zK�_��Mh�ĕY�g�9͙�p���&X�m�S�I�	.�����5���6�Z���q��lw�=is7:� ���ɺ������6֭h|D��H^iBI>�)|���:���i����Lw����n~>���d�]��Y��S�r�6�P�oY7^LaL�$��r2]c,���S��(`=����c���1~�S>��K,�b��]N�5�SD��u]�T AvcM���4�a!�/��.�-��q���Rg��Q�q�]�(���U��d�f���(�c?��n�7[�4����ϯ���_���e���{��ykM9��z���Z�o.Z�a����ر]Ξ�}S�y�U�\	�4�~FڔG��"eȇ�������$��uYIX��>&�;2�ff��L�u��`~ą'"P�!R�s�4XS��UZZ�l9KX7Q����)o�=�l���Ԟ��gn��K�g[���(415�N��E���z�JKX/	�D�k��g�*#_��r*�0�W���x����ag6]���oy A���3:�7����k�d�f8�Ђ#"�],��%y �>C�jwSf%��z�Җ�nY>��<�j"y�o�o5;g��IG���g4�hQG��uۄ�� >!Em�r%ZX^Ŕ{S6�:�.m�ofK��Ͳ�[o����n��ڰ�����<��{���V���
\4M9��8�h�C����I�&�OO�l����7w\2J�9])��N=��q��jP�;q�q=�7Ų"a�����P�\��ěK�;09~O�V�O��p��Q\\O���.dw�'�Y$|�Wu�&��x[>�Q�?�J��T/��c��a�u cd�����t.q�N��=��8�%�N\����;�O���a�O!��7�HSa�IE������P���{U��;/��"��yM'�	v֐O�r�t:�����P9�۝=v�cY����X�*�+��L%�z�Ü�Ͽ��������Z��<����E}V`1OY���ik28���F���H��\?]����YZK7!�|*����f5e��ڻ�E/��a��ryh�����Zt,_�ś���D�����L�w�'��WH4J�+�kr�]����@���cO�&�צ��u�(�/���k�Alt3���ЋL�A�5
�)j`�]wE�JUt��G�jp�H|a�L�y]qs5{�\#���Q��Q��G�#jw��'�}�������|��3��I:,#��+�>k/���'k�PV%�r� U�v��T����q�+?'t���4 �g<�� �(v�9���G����CW�r`�7��:-+�ҧu�Α��U��T���9�ٌ�G������������#�(��=U_�O����'�'_�*�����nF��1k��%�%�Pq?�xzc	Ũ���f��M	KT�j��?����T�)7v��l�6W��=�����q���M{ ���a�qI=p@gq M�m]�5jN'���Lᬏ�ݧ*��9[t!.]ܦ����96�X�����[�m����R����|o�`��lB�2���N�ǋ�Mg4Z1�#�K��BEz��\]��&�Et�T��,p�"�	���/�.�*����)m��`�����H4��U2k�F
�:{�oo_V�F�{D*M�N�>�gI��oT4hoѳ�f���Y��!�hz6��ŀW{A�0�:З��q�t�1
��yk��֣d��*�3 �hM�QA�"sDL<睱�ݿ�R��U��.��=���z�Ƣ�G(�l���I�ya�l|����b��fn�x�B�$�N=�qx{��|��m�:PTh{�&;9���l�:ʘ��1Mot�f6~d��|ŧ��^Ҷ�Ifm��q��khSv��=���\�&?y�H̠��(�6���b	$Su�^��=B�_"�Yl�l@@�j+���� _���'K3{�����B�b*������ j�;��T�#R�&V�Bq�)����\a�����=�m^
I�� ��o�8��E�PԖ}`�ʒp�����_*Sz�҃o��̼z�@{�E鷧��r��$뺣��&�i夣×�<��B,� ���	g7zGf�G���~;0��k͢HT�F
��o��<o�.���Ɩp���Y���0Z�B��z^�g���f����@w|R��0���Մ�r�T�D������H���'��1{E�����	��'�e�:CD6x�$�HgJ���u���Ĭ"!���\�Z{�� ��Ap苹8T�T�v���_�1�&��7��c��A�ݝ��Ӗ�qN�Ē2�X<��9����<��Q$}�0g w��z�.'�ž��C.��	$8YƢ.�m�>���\q(���kZ�g7�4�(}������s��|?��:u�G2��)�'c�u�i�۝�Gz�ma� e�JN���sa%��h���p��jhM�m(V�.�����b�a�o���O�B],�(c����U�L�4�m�H���o�Q3���8�ʫ��_|��N�?�	��<��#4��Lգ=����R�w�P��Iw��A��}�
�]�o��2���d�ǀ�*o逝�/7*J��� �� ������<����{X�i@�!��k�tm�2�B��#s�ON�%����ώ|GP��U�_��"�F�1.�xB23�t8�E�G�ו5��&�Wx�'��:Ca�@
{҃;:lPbB��Թ�A�n'<�$nIB���D��C�l�V)�Ocld�Oci�*-Q?E��C�����{�@-e��7�c�i�&9�)� jH�`�2'|ϺD`�� =D	�Yɯ����^Xi8����H5Px�K�@TE��e�4��./A#��8��'Z܃
c<p�������ʹn�� 2+�ٟ�_�+���?�g���>�.�����)�؉)��y�}�H�X�?��c�T�M��ѣ��y�A��Ű��Θ�CF��������ӻ��t��м>X$o0_����!��1d���@�* '�\�b��(J>c�m����������D�Y.ƶy/��-VkN��Js�6<%E�2�'Џ����E�����	��8�B��� ���z q�L�Ă������BƤ+�y�[�+x��T�b�L�(",�CDV�$ǵ:�ꇌ?��@g'��BE�H)}s�(���<@�pc:�FVr��u�9����*!��w���fA�v~�@o�(GC^�hn���a$���NF�+"�O�"iJ��uK����}�.�ZU���y3��˩c��2E ��Q�Ք��>R>oȧ�7�[���`0>#�+
���'F�/�a�h�����J��L:���\W*� �׋C�U�T�`����k��̼1�W�ņV�.�����*�;���bٸ[�|���D�"r�dZb��ޤ �����~Ii����>�A���.Wg���J����iQ?擄cp��������\�gc�19u0��J�P�`ϲp���X^f�Gs6Q(Q��{M8���d��L��w�i���9�˝nϠ��=&m1��>�§�\d-�a����3�ș��\��l3�$�Q:�Ń�kX���<���w�1�T,۸+��b�S�Ճu��V�� b�����՞F��s����cb�=��ڥ�f���ʉ<���L/WJ�C���L9�0��7M�9sh�[���[\�+��2��{W�?�F�v�X"	,�$@QP�*��PL��~y ���E�9
(��e���`9A�B��r#ڋ��T�zko�bB�5>YAO)�~��������[=�#~�
�p,٠�I$���k�����	�G�n!I�J��Cg�a����c��iT���)�Y���漭m��m}u�����¦�x"4\�u�B�H���-�X�3��y�a�_Ľ����UM���Q��K@�y&jl�6[
; ���tH��i���6ῷf��g�s������g2�p]9����|���G�F�j K��9�Y�.���;@{��yVA��5ܰc�H�n��		�W�zU��c�7q�z{2��Ԇ�����O��i_���0�?f:g�J��m��Q���_\���2� ��Xy���,4����9�ܑxgz�ʹ�>�>�>���eW���E��)k�1>_�t�v��M5�aW�K��πK�k9��ߎr�+��.��kE���rpU���J��=��i�O2���ӟ�5�_tUx�]����O�wD����� ����l{8�\�����6#�p,��	=�����{���O�i�;�x�%Pt;�T}�K��al����"�	5����:t��pͱ����[���GY�<����"�����#B�EI"*җ풜�.�V5����R�����2�{�{
N�k,��Vs�T��Գ/!�Xj�9��N��JZ��*�/�y��O+�l`M�Իf�*�I��2nB�����CCaK�؆4������z��.���b�ts�\����![e�e�����/	�����D���D�z�ВZ_��9��lڬi	+y�*�g����>2ɤ}a/��N\�-=/��N����r`XN�$�|"����E�K�㿽 �/�
�ST7Io2�t x'����[��d?�j�]<���i�7*��Hf�&hUd�Q�v1/�MBr�35���6#�ӼdI���ӥ���(�|�_��b����띞,{c�{�OFZ@��R�7I���y��7�}�������c�0�KB���F4a�Bn�bC�HD�Z�Jv`I�<���r%�TW��Au�ed�k�63��|�Rlt���2,��S��q$���>w.��{��O�OkÑǒ�݁t�Y&I�_ &}��
��aJ� ����T8��u4B�ضh� ÿ��Cx;�����/���`n�G����%����M���[Y�i=ԥ���������r�xl��6�0��������p��ǎ�[���DT�u����:?w�uY��*2Ǡ�te��H��"*�
�`9�4.T�ŋl(	]EI�g-��0��"�����v���kVv��9�&��ۛ8
�1%'TK��U�Ha��TȽ)N�֋\I{ӑo�7AX��1�(�NB~īj��R�%`mt��Z�}���0�ou/G��Z���l�]�`ٯB�Nk�Tڧ�����������2�8Nf�
��*�G��oZ��R�[OH�N���О,()��k�Ԝ�e����hIZU8�)�	���^PK[��'� @��xi���L@KZu]��9�BX���a��8�@�j��U����d`�F7E�ܛ���nq8���<�Å֙>���_8¬�L{�[m�hڰK1لV�wO^xkZ�O�1F}�ʓ� ��[�m�A@�K����X�|.tE�r|�o-Ϝ��f$���y�~#�ވ�T"�K�)�ڧo0M0��Ό��͕NC�~�U~6GM��-9���҆�?��" �$�D���n��������`]DPΐ��(��8#���
"�Ѯ�:rą	��o�8B��]���:�ތ������W�Z"Y귳�ߌh��J^8M��)��N�8���r�Y�MH�>My+&^���pe��3���:��TaԻ�-=���Bqn�׳��)����0۰�����y[��d7���v)��]���2��F:+p��8��x*D��\�4���
c�����G#?���M��pھ��kϐI��s��].�n�1�k��M�,�_�n1Mߧ���·�d�e"����{�M.ɞ���Uǋ.��X�	���W
ǘ�,Ӭ�jF%����3�Љ
j���F0�kX��r&(u�qJI( �-��ٞ�J3~M,ذb�@��������!��H��t}I��7Iգ�4"��(�e�˲�+0�_�e�K`C躪Ȩ��N�<"X�������A��˲3M@=����E�Ya�z��� ��s����X2�T@�GM=�ƞ�h�&cD|�-�85�d\*���4�AĊw�:E~Z���3���5`�>���ȣ���E�迅��(�Xױ|�
:�(�`��&��V�;������!3&������9�f�U��F2���A��J�"��g1j)��d4�Y,�?.����^$ّ33��S�`8f��̶/�B����Tt��HTΚ��vw�Ⓑffb� f!<�+�u����6`��Qr4DR3K&Xg*�C=8��vp��[�y˃kj���sa����/�ҿ�Uv� �gnj��f*��Y2� cR�[��A�.�	��>�ƥ�!b�^���Y�L�;?dĔ�?��.�`|�9R\{-\��0�R Ĳ_���Ei;���fW3q���K��r.���p&�c[e��OЏ��⶜;ku�,~��L���,����m�:�^'�V��Mz͉$�n�<JK��a�?�b`� ��+��j.��q[����>�}�/��>�g��p-���AIj*`�g�!���w�ق��h�o���i��rmA�y��Y���R�E���+���o�ƄL��������������:�̛�L>y�.<�^� Sy���\i���LeR�P�̂���v�k�l鷩~�k��5������(���+��R�	�\se���/�ʟ�xVYȖ�m&n$>㏗>'Ä��Ǩ_���y���˭���UR�^�;�R��8!�)^G�C�*��ȓ�P�����t��:Fj\�5����	�J�RV@GJ�"�qF=�$�9,yX��FW}Ќ�(���2"�34PP1�#�a��Xݪ^/@���d3��9^��u��!髩ҞڦZʯCK�p�?��Mr$�I�k�����u�&���A#�tܨ�,N�x4�L|N$H|��H���
S'�$�ߠ�lA-��(m�<գb�������IKvqL)юF	����K��P�Z���NyT�zuWO"	�(1`�ۿ��s������G�=,{-�]�C0�D=�@���XN�\���>X�Ȣ/��(ݯt�.�ƎGhv��m�s�S��Y�a�Σ�����?�l�
��^�����8:�C�8PO�y?�y��̨���Zfs���;�⡜K�[2���/T��77���;��۬S���Y|�>a���#%.�lq������i@�aЪ"��f$g��V/"դW$t�������R}d�'�&��]��o5�}披��сM�E��v޲�)�d#WL��Ե����DN��uLO�D�^j�T�t���ބ���swZKΉ���Vd�4="ޙ�0`�\�n�fs�A���tO�G	����J��4�a�>+9�ŤLNA��ގ�-O}��~�+������g�-'�ҁ�����ȁ5t�7��T31�Vh����Oh�,t	4�q�/ ���(��	|w��&�Z����~��%�������]F�ۅ��t��� �"���I��2���O���,��`'����"�F�/ϔ��F,]��Xdm�:P�C����;�g��*�/6@�S��9�t�p�v]џ1eu�~@���T�T��#s�wʂ}����CH���q"�3��נ�ɱ��Y֘bQ{�ʅ+��\�X}�.���u��M}��NvÉ=�˚��\CTE*`�c�#S�ܨ����Ac^��ఒ)>�u"��)��4~��n�$mu��E�6JucL�z�Q�
�����'
������u֧�|�ߕr���EY	��{�]M��Pg����?ĉ.S|�a��R(�#㜨�у�j�`OqO�	֫_K�Ч�kv5k�ϳ����7R3+��)��XHf D*��E��n��FCP�t�<�E��w��=���Q,��0u����?s!-n�������%C|��3�Ic�4~��7��񜊑�N|����ťϺ[�S�#����q�����F�LC%�����w�pN�]v�p�-c�avt�,J�3nӑB�1\�?1?y�z|�	~!���Ļ{��\J�9�T��Qf+��Y�WPKSc��SE�<�$��Ժ\�C��N�>%�Ѱ�[cUE�c\6%�$��KP��$���(,���ǖ���T�����2C��Ҋe���4�g��Y�� �U�rj��Pk�8�I��Ұ����,����#T,��X)����k��*vm�ͧ9�L��[��zԁe�e0�ԝ�|.��	�.;�����T��gn�<���_���L��l���Z&>Fwu"޲ib�T��l!oZu�R%JK�I~A�	Qq8��ѹ���Ⲷ��!�ƿ	.ڡ�C5�w�*H�D��6�(!o[����V-���O�V�jx�pY�K?$Xd)��-h$[��N:/=+u1�m�~/G�۲��:�J9�����̙\�?�b����F�f�
�8�O+��A_��!g���Ծb����P$y�7Rx��j�Z��?mv�[��vVߒ�!%�R���q�*�*;�	eJ�� �̳܆~F���E��>Zsl	8+�y��f��~ϖ���RѮ0onv�x��%��ne�/q��� $��v��������~���S��N�8�tڅ�0�z�x
�o�VPxx���Z�l����m'ji�r�Ź% ����}.�h�C��$+�=��ʡEp0�
z���Y�$U3�g���xe�N)��|�B�� ��{#v����O�n����+��R��~N�|��;c >%���<G�������{R��I���<���DŔ�\#�}稉ȡ��Oi�P�w(d��峘v�×����pA<�<�$V�6{+��ԝN"��&��y9����8������J������ɦ���]̔Y����`Ƥ�'ʫ!M�ߌ�����G���o��>��"�w^ߣ�,rc@�͞O�]�� ��5�z���,{�5¹16?G�n�wg�Tm� M�A���h�*Έ����R��O7X��/��h��~H�su����\���]����*�ef��M�qI&����O�^��7[Bڿx�����hߛ�~���F����y*�h�\�G�3�קvk1��,/�A�9�a�����!ũH����H���!�_� z>K{n�Y�FE"�1K�ɭi<�nZ�b,~��>�l�|A��='���[Ln����W�>;���*5��`����C�k�&�w��m�`�e�";і�f����/��.r�B��DU�t� �wZr��go�j�d/ab�.C�S3��nb'���������Qd&�=�veI��Hi���̉��3�9_k�8�����2�u��Z�7J���!�3�����#�A[� }}��ؐb��*�-�����qkE�0y�����ʉ�-��x�b��fo�Q�e��V���$e�?Dv�gwb��|V�/D�1/�s���'ބ�@��YM9�)$|�����s={�4uc�P�~�ʗ1���S�<`c��*O�S��Bc�N��A쐰�5J�8c$4�y#���:��l��)�=6�4ª�>��p"?Y0?�s��X�(NX�@��b�$�S4�u%mL�I\ҞpViZ�0p���X9�V��m��Ak��O��d=�;���u���c�X�*���T�qkBPs�٢X�ῊΑm���ר�H�qՁĀU����2����I+��{.�X��*�������&�,WA���6E�j��O ��S��O��ߋ��C��y.�֏��"�hg��)�	
@ߝ#O��}���"�>���|o��YT�{9�F�ָQ}F&�,yς$��{C�_�e�P����g
&@��b�9v��ISЬb&P�l�/@ݤ9�|�����ʂ��e�#z��a�|��T俒A�b[�.�ʶ�R=�?��p�o+�!����@urc�C�c�\j��]��ۿ7�@w�?ʊc��]
���%�?Xd�a��D�v�,�!�:����ұ�ٻJ	�7�ں�i⋂�����$��w��R�I�l��X��(Q�ô ��1���Zg�~���Ez��I)}�n��$O�_��<�{�W~Wl��y���� �U�H�����F-
�:�Z|y����A`3u���x������S|�0���̖ތ��_����?�q�`�
��aG?3���i����㊷VY�����υ�=�S�cx�Q�u�)@0P��:�/V�b����|[�7��6;�s�I&,�ڧ�8��n�t�;�kαS0*����d��������~U�7�7�RKvD�$5��+�_��#88^�ED0�G�N��������'s�x��˭SmN�\v�7�l�6��'9����5wf�)�ב�Í��A\��.���t�PF�XZ1f{�f��Ӟ˂�T
�ߑA�$���sĤ���7��O�H�u~���l�w�!& vHz����)�bT@�\S���7�U�붪L��B�jF�[c�Q
uD#��gGW������-p���Jy�k��#��˙��}�t��8��w/�J ������<��:�q�s���z�ɀ0�g�	����ۭs^����~G.����!4�֐)��7zS��·�|�
�.Gw�d�)��9��ƾ7�٘��[���0N8/�]t���Do�Ԅ�Y���^�����"fAB�K=��T{y�bm�_���]�M��E�����A�N>�گ��>nd[Ǚޢ���=k��0IQ��B��!��̝�7(�Z=2��[�|�}j�':f����|Q.�nD�:�Di��@��Q�&�J#�"0i���^��+9�z�ƣAz�������g;̢��w�2x�z85�%�y�N�[����
ͳ�Z#�O��@xQ���R{ z���M���h�B��s�����OG@��m#M�m��&5����訟|`�N
�	�9�L��+\�O��dD[5�˄l��P�&g����z�=d?@�믆c|�jzg����C�ċ5ζ1p�PO�����yPx�5�����ӭ��B��K�-�ɗ[��3�AI_fB�6��QJ�4�9�F�T�V_�%�"�IO^� �0/A� 1ȋ�ۣ���>9%Vn������M�l��̭��1��Y}o:�O�6�E�Y���"3e�C�`�7w��%u���e��&�Q�꬚z3���4� ��Q�{�����B�t��UsL���V}�o���9�6$d/U��T^���A8�b����S6H1u�Xqk�$���j+�R�qu?ru��#�Ĉ.�r51~!����T�����e/�)�ۀ��y��c��QX;x�Z��R��W���<	�&� ���?+(�XRr~k#�T,Ml}b5�[Z��]�kĭ_4��⃷�ic��J���V�尢�#YL�~c�U���)BG���O��96�U.�t-?Sa��1�0��7ցa��Jo|J�BItα�?&�muxP��z�� u���F����s�N-2(�m�܊+M�hjb�zo1fK�[ m�rB\A��� �2�ZZCR�ꙴ%9Fl��[O�mw4������C7%�Z�����l�@M[?�������5�G'�:��bC|[_+k���^z����:���Pu�Mb�ơ1�b%�wk�Rf�Rw�y��>�m�?"o�ªE�T%c$���Pq���C�/�P}���{L�}�ٛ�(��o�O<�{|j_�t	�揓��@��@d�Is֕\�q�r���KT�V]�HZK��Λ�\}�7Z�A��������B�2�h��� ��T��m����Et�Ѯ�PZ��j���*�`
�Q�4�J+pD���6�Q�~�3S\��TY[/���9M���^���r�?���Q����Z�nʂW��1ʦw���	.5?c76�L�=�r����^u���Bu9%���J��Ա����{	����J��o@����V��U��$+�B����.�h��g��!�yJ8.�`���5��c���_�����w�ɰ{�\'A��xO��3�NV��*���cH5�t(�V�����R�Pӕ���]s�~�U��������8��Ok6��46`��J&�nض�nx'_�I��5���w<���?2[��CXޓbM�s� �>+2v�����t�_2Ag�'5r�\��ɬ��xkFL�&��[8�q)�FdG5=��� �#t�a�0���^�ZxjZ)���/�x����>A6�R��ؒ�I+"����3�Xl�v��5W����'�]z>,.Q�ݖ��9˕�_|\���&�'�����W~*�2{�G���A�)��~�ik��+�Zٻ��H��J�$��W����7�d� x;E����F)��Z���*A9���D������p:"L���).6�75�9�;B�ޞ����M�2��ø�G57�{ne ���~��UR|�gJ$IQ��ͥ�.sR�x1��s�s��Y
��8ȑv�<3��ry��Pը�u�2"��Q2F�, �^�`���^�
UE9�B�zm� ��P��aG����2j������Z�'������)˰��O���Kh"���'�P��L{ߕ�������c5y{{7P 1z��~�Y�R����q�9����]6x���Â?w����xX�кխc���~��� �% �!,l��4zͭ������?)yru�9�K��v���=F̶+�J�GLg��>������7A뀩?z������k=����SZ(�`s%�;��)#O:���lI������y�q��Хy���gU��"̑뺚�M�_S�20�
L���0���&ܗ�Q�k҆D�{]J��Uy^�L���g`��m��gvMR��W)��@�ܱ�w��N�֜Q�Y���p�9N&&Ǳz��(r���b����zRds�P肥!a���
���k�
�#��/y�n��%s��7�!�+1Z��3�z�~�0[=/�XNg�ʙ!�C�ܪ��&�A�g�	���C@} ��#X��sI�4��a�����[hW?�_ (�g��Ps��w��ܜ^��0V5�j�#�!S ����j��!��[wX�bD+��[���C,H����jB��/E)�/hL���(�]wʴ���a�en�5RѶmt�O�� g���c��J���2fc#��p�k�<D-?Ǒ!�sMf厗��gq��8�X.��7�����i���gMO�Qk3������e����,׺rV!�Ⱥj�&�>1N���˷k��A�y��:�q�K����E��.�/�%�Y#Jt-�Va���;n!�n߯��XjX�����(������6Bv��U�<��<�M�t�,ѧ}C���x��3�]�#_���+:�V1"��j��)�s�/����Y8�V��z6�޻��u�I}������V�{��w�Z����Ѳ��$Kw�p3���5 %K`ͦ؇�"IBߒ�����l�lF\�O֊�)��IE�a��<Np=U��m4��c��z^[�>�BN'��F�/7h!��e |���1�%��֤��7���w)�ҙ�z����S\[�\�-�� �P�B&.��|8�Rg	��[���޳�Gۂ=�s��1R���a�~{�S��I��x&&�I��I-�\�F�%��a�L;���9�{	ҼJ.?	y���	1�	>^z�o9!�'B�,7HihsA������o�S�`��,�c�zh7�5{�
Z�k���? �gK,/=�`��,�n�\xlՓi��c�T��lC*���"4�����(Ԫ}T7t�v˃w�E:���*/6������I��46O�׌�����y��J������#���M�[�J+�k&��oQ+��o^8��K8��
 ?&B|��l{
�J�Q�a����8Q��s)LEb�q?����~ś���ϡ`E5���ǐ����3=�
���e3�9E9��A�
�,l��Ԭ�i�!�(*-l�:='B�y�hV.l��m!m��,���^�e|����O�,$��W���Jwa�vUT~�*{��A�6D���҈���q�X^+���5QA��(+�J�a��l9��8�|b^��_A�����'��m2�i-`���"=��_������,-1^MYC�����ɽ��k
}�u�%�!^��$)n����[��n`��2�p���Q�=��?a�\07�z��L�;]�Kq��:��#Xp�x^�A�݀����>����ȍ�����:Ƙ�����4���cV�h1� C0n�BB��k�>?��c���F��^s�����_�����1.�п�ķ�Q�  t�d2{�N�0$Oo����j�?���K��#g�>f}O���+�G=Yk�=--��gO>��M��C��5�kCɚ��8�v`�_�����_��3��K��/�l"�4ό�����S"V�0�ݳ�� �1"��GO�)�_  �n��Eۗ�N��L��4�����i��������s�6�n��._r������M��
�����r�w6�t4�Nf�冉z���n @7��%e��X�_֋�'R֯���2Z�UlC�V����LAm���%l�}_��[QKO���7�,"�~�7��)��w�(�s�d�xh,Tΐ��Wڄ~T�BJ�Oz�E5��/߿�sk�B����쪆��� ��`�3� �c�5�U�Tɀ�r���o��d%����YcC�.�V�l��θ'<��=Y��o��q6g� ���H��7_��UA��%�VN�%�6�g����ޣ�֮�_{['(�[�zϚq?<�;>2&xU��C1M��g-���b�PB��E�߀��`���c�4!S�F/���:ALd�9���i�L4q��&��S~���J��.�[�f�m�2N�sS���<[%�p��1D�X�ì�����?!0m�!G.K�.��DK+�X�L����ݥx�֒eӾ�e�јֲ�(�`�������&b:k��1/�0΋й��'*� %��/rX�e�Bn&~g�~�.!��
��B#�˩-��.<A0���^��Q�{��u�m&C���G��I�[P@XU�GO~��l-W,cI;)c�<�#�����?�-�"^�����ki���Hd�?�l��T�*.p�wf}�6�1���� �FBy�i$���Hn�Ey]C���!cZy]<d�[ǉU�i��`�"x~�ϙ�s�a�w����}����(`���1����8:��5	�	�hf��(��uu9P�y�v7����k���XT��x����@\�iFX��͎pSLXW�6�ch3�g?@��C��$�VB��D����G6 �RbksZ�yėH�qh��O�p=�:�o,9z�>���l���:?��'h��oE�|%h�&�!���ϵ��,�W'�>��|���ԢWo��J���Dv�(T���t��i��]�4g��?yV��fV�q�W�6^��p2)�}��dWM-5 ��������au�ࡄ��_ˑ����V�1���t$�I��o���u�	��/�P�9!7l�E1��6o~�%ٜq�٥=���Kr���As�W���9����?�2��"��MC��R�ngX�
e���ʕo͌&&�uG?�S_LKî�cg�쟍���B�q�%���'m2���`��G�i��nfRe�S,���W��4)=�(�׉V���z����ߡպ#�p���n�`�Y���M�3�:�m���p�
�����C'���9���g:�A����8�O���D^m�,Ct��3�m�N	��D�=�5�#���ф�D� z�	jC���$�o	潇��k�.N{�W�~���K7����$N�3��%ݒ�)K�b_��+r�B�۽�Ş`&B7����y	i�(U�1!ؤZvwm�[M2cg�&,g��s�/{LR� }����F&/f������y�W@������/f�_��u�N�;��� Z?3
��Sr��t@��	��"U�Ϥkjx�e;���"G���G�B�{v���ֵU(&a�b6Й���0���|ƭz��zq�BOiعrm�Sb�v�Wj�5���x�a��j;MCj�Ӓ�o���Y���s�CO y��-�{�D��P��We��\���X6E�2���;_DLf$�c��Jd�Zv��^�ïj�g�?�D�2S�'�ț�`��q� iZ]������A�����󀗶���!�}W��3�������N�P�d�0� ��bf�*շhR�����+�ߠ�2�(��MXЪ�5�?������Ρ�^��BV����	0�����82T"��FwY}�j6w���G�+�Ǡ��j�n:!S����ma�o��WEHS8;��|[P�,ū���w��%��,{o2��*ԣ�����^���e� ���6���|x��17%fȫ�k��ґ�r�Fbk�\L�j�M��3Dp�<\�޴<e�!Ի�3s�1��?�����<we��O�)�o�!��f�Vx-e+��b�����]C+�"��v��O���ֈ��:ӿ�&?ey������cA��]�&ȕ|�3N��3�X�r�-���� ��[���Q�\��q�I�5ټ)C>a9}P������1����"� ��s
���m�ŜؠM��~��c�N��c`
�����`�r#���j�t,�㪔��o�T�=nz�9t�W*A��X�����g���eܜ�����V5�3��s�TysPL���B���`@

F��Y�B���c��
��]�*����'"�>K�	���f��Iy�Tv���
���\~��_�[��Y4���Ew�����{;8��9BS����%j���l�ʪ��#q%m7�q���8�K�r�$���<8~6�lwdW���*�{�B���ꔨ���)�u�c�����*����ڑ�g�8%u��:+
�{gB�'J�L`/�/�s��/Gl�i�e��B��Oܼ���P�Ųl��%��z�m;���vR��Aė�2x�(��o�
7�nZ:��F����vg��N P��^�j���[�������T��7H���:Ed���ϩC�T�3܃��JX������}�b��R����9����0�/w�m�@�Q��8�$�lIY���HY�����E���l1&'�O]k��セ��	��9����W�?��T	Y� ֍� ��^�>��}��Z�%>�
�:	��*#�urC�ƈn���@�[�6z��;i��.R���4iEa���������+�䌺���gi�%�
l�3�O)H��S�������&6Y"4va�3�f)�W�������= nә��u�}=kU8@���T %i�_�ZJ��"�J��pB
��o�.J�@2ߘ�)o��͆�Vo1���� �bGग़��U�	rNL�8�VG���}���O.��=���Y�,#����
~sA����d���&,��8��=W5�î`g�]�0��L h,��H�۩X���/�mr��#����:pi<}`��9�v��T�_*|���	�DI�[�,*��o��<C���Q�{���!� ��BS,���B�k ���1�n�l{��lQr��
l���s(o*P������g�'�]���kp`F4~^�E�t��޿�	�kA�<�{t�{6�f�b���ĵ�Gf���	rU����gh���3�Ҽ����>��-S��C���Ut���4l����,��\Xy�-1�3�l�D����o)�`�A:~&��N-��׾h�25e�Wh�^��+I�X�n�@C�Eh�l�&��UKaš�o!��t�zZ�,� ����n�e���E�!T��R#/�P�4W���l*�T��g}M�T5̳c�~~Q���&�QsB\C�]tM�Kk˂ߣl��:(�FKz���y*b}fz����t�^{�}�h]GЯ5]��ۘ���i�O:��f���-g5� h�j0�����L�1�JU���V▄���I�d�B�w���Af@().����Q\��_�C�F� kהd�J����΢ǖ@�<8K�y׼�p�y��&���v�S�j~�6B����sj3%d��c�2�&��GRX����#6.�{Y[��t ����Q�B~l��Lz �e�po�Kn�&.���B'v�tG��TU�u����Q��4Y�<mhcpj;j���4�Z�,6\l�" rm�)#�ټ��~�*I�-o�(�L��x���Q1IS����7��-�yѦ�SG�1P9���Ry�|���m����(�X1��0Q�9�p���e
�s?lz;}V���ӥ��SL<u(L��J���m�xu�juП�W�{�fo��������TRف�˱�V�֠A�"jd�ɇ[�kG$&�~��� 9|�͡aRU���-�����C�C��(lVz����[,�W�R���_H��.�B`�u.�G�2����O�fT�q��H	�23'8M�������X�Nm7hk�|���^f�ћ�;��*B�;�xt�ʮ���!�.���iS,�� �=��R�7.P+�H�گ�0jk*t�27�X��/���AB�T���ȹ�/���@��Ō���~�Xk�=�P*�1��ҳ�Z	�H���@���`��I+��nD��L�[~�qE��#�Ꞛ#���tSW*_���j�r����N{���{\�[���s��W0'��)	A
����C`�P�彝���0~���'�`<��kl@���x�Jf1k����F�d !��ڰ/3#�^K�,7�ޔ,��r�s����}�Y�LŁ*�}X&��I�c�>ݳ�Ӑz�r7+�=�Պ���B#��`�V����? �9��|�5���q���A��)o��-@��C����`�,����@��|����tq�V�h(M�+�9���?��4�q��	˴�	�'�=Iz�u>�[�GUQ�Q���[Avo�բ?4<M�/B0w1���Ͻ���"F�O}�a2>���C!���.B^���SKس�E����7�
$�3��k��L~ضdp:fp
!�� �iƶ�F]�bS�M�(���:��j�&���N�ѸB��&��F>{��oOsIK���x��2
SU+��J<CĴ/rk�~)����;k3k��_�9+r�h��!vQ;�kh��u�p�Q�o/t��:��z��%�%���P�iBC�����t1\����1��Q	�Pi�fOR��И:sv��eY�im��3O~)z~��)�Ҷ����X�QK��Rf�(0����J\z�;��vΞ[ z����t�ۜ��r𣽆4t��������2./����,���'�o*����%�ݽz⏀���г� �Ȗ&3LY����D�K��0l쾔8���.��ӗ�]�T��;���&R�7t�.��,N��ւȀ���W�`@s��R'��%ڜ���݉�Xb]+�Yl�K�	�����d4	�N|��4ӽsMt��8f\	2�WS�p��6%�l�9sƆa1%�N�jM�&�d�o�B���a�(�.���;'Sw
�EW&�V�M�Qq���U�� -��;�mr�;�Υ�m��[=f^�F��>�wr~�(�n����pA���jzt���
��~�,KiH�HW�V��`,R[����#'s<��RdDrM�(�7��������C�3F&�K���؋t��p��g�+���P�����7?���\�`�;�6����Vu03��~B=���@�g_q#ZKE��7-�����& ��m='w�=�p.UV�����!76-�U�W�zX�YF/N�}����=��ە]x&�P�x��fM+�!���z�@�V��%�K�f\��&�����|��,TK�"bj�����Z��D�Xx�%��$I����xAnF�E�)�÷p�K#"���e�i4�Ëy��[�\^+�΋e�D�=n�#'T�}�γ��+R��z��9��'�xɊ�Bk\�Ϣ�����*ͧA��PP�O����q��!ث�ÝP7t���F�j!��L�i�:�[�C(�4Z��i�oƅ��v�t������4�Ҧ� �Hǝ%���h@� ~?T`NΦ�E	�)��)[F9�< W-�c��@�u&��=j�ljﺔ����V%�9��BF��XG��yd�W���_N��U�s7�P��nh���$����LY=��l����Q9@~n�Q/���@&��v]FL���D���y��
�]�@��{�[\Dfg*�z�,�*�S|E�*!��J	d{�����M�D��BVj4O�2w��VL���J���T�!��B2Ɖ��U��5�:�Do���}I���}I�o��f���#�G��y@�瑮���_:�JI�Q�9E��y�H>Z-�� H�cӋ��@�ٖ4�ʊ�e b�k��Y��W��<����;��&	����"C��_������<�����Хh<�1W���}�A �ǘ�j#�)
́�����?��:8�R?,X�m��J�"�`|F�T�Nm�/�7k��xʧ�e�G����YIw�*����տ
f\#o���KA6n�FO�cs�*�L΂�&9�B�i6�ܖ��C�I���\��`nh���!���o�$��(@ק�Q�{Z�83	N�y��Saoith��'���n�\���ex&!�ȣ1�20�Q���4c����v̡���<I:����ƣ	�+�M���(�`�W/�w
u����� ��h�=���r���5���ؓH(�"�l��I�_v��o��"<FA^Z�K,���� �G���Y�ۧ�S��� ����_�uT�&L� ˡo'T����[�ߴ���4þ��{�Ȉ����A���V��=!�K���Ag�^� >?8dF%�"��^,��7��*1�j	����p��ݠ<LS|2����аB��O�6�m�[f�ms܎��	��dC��V��7 !o��K��ժ�`��FY|�a��Cr��$�|�y���Ja^�;�)��$�# �"b4����P��W��OԪ
��R�.4�K/��q�~��oLql˧���OOK��ǛB]M�W��SjXlR��0Mtg�����ۊ�Ǫ2P"6۩v[%v��h���``s�a�=�NP���t|�aޤ��b4)�O�z�G����������y����[W���V�m�T=�xJ� g��] ��]��Z_����r�Ļ�Zp���f�4���U�����CH�e*u\� �4��i�9փ����Mu��[����&rKJ��
��g�%� �4ɶ��zh�n�q�:���P�,�Ը?�2z��v�X�"
*,�����>�2��E���ͤ��vA����YG���<���F�}i�ʊ�'���-�~s���$I����{�Z�H�UvC:d�O6���)O�&x�l2���"�m^O��*�d��v�-�G�3����G�xi���#����~��<���f,M��֍7�!B
6�i%pv�M9���t��P8{EkTE�f���[�*�q��1�'���!��7��K�ڸ'�JG���=��Iv�Q��G��p']�tԼ���0����G9��1�hP���õ��$o�����\F�Mx��S��4ڀ�k���!��O�r���V_Y�]w��7��F@��C���~=�{�Lų<�/��AG�=e��dŊV�SsGw�PziC�����C��C���J1H�A���y���P����>�WFH�ﾌF��F\��d�$B�ۋ�aq>�H��Yi��j���� �Y�%cTq��"\��4�y ����8lk��j�+�g��ֱX*?��`�[/���ꍖ����^7��a��H_f���0���[WV/����L�@���3�A�R��V��DHI��܋DWƈW!b�����U���z�Y;V<�]���́��܆Ŭ�ȭ^1���T�eD�*��[�#�9gt����ZӐ��7?��\�I�N�� i���?���hX�໙��e[Y�u��dN,��!=������]�1�R�J�T�u��E ;C��14��$�͢����c�0������!#Or������!5�gDv�*rt�ČPY���lF�B8B,f����=�/vA	C�Մ�=�
g{1�'�uf3��������>��/��rL��^f�@CJ����s�F]T2�/s�R�Uz`�S����:#��Q��͙�%�U[��	D��odɩ���p�: �v���{BJ���2�*��l�upZ*�ז���]�	��02 `��\���5��&C[�k�4Q���Gu�Ц�!����3��[\������Y�݈�@�]յ�0`�ʺi���O\D���M?�T.���fh�����_R�T���K��?E��nb�?���=�2���ٝ~'GU-���V�lAN��¹�à5�c�Z��.��3�$w
��G?Ӛ>ZW�2���L��k�{
'�,����(Q�R4�Z�I����[h\��S� `q�Tv�R����8/��yO|��sAh� E�����.1C�{C{��r03��e$I��!�i������@8��Id�w.jN:yn��.��_cm��;T#��1��F-�p��{GK�n*d6���G��Uɍo�E?Xһ
�1U=au|f��<�}g��*�H�S�\;i�9�p�#�W� ߷ÃI�-�Cy���HK�y��'z����7;o�l�O���<l�;��p�T��N�>�XL���������d��$�S�,Ҕ��x�}��(�>����Vp���f"K$�Q:S3��/p3��<ԿAm`�+����|lK�;,��(�n�8�G����������sv��J�SX
TVN����q��4!s x�X~n�-P���j"]CTf���/�NIM�_�������lK�Q5z�nM,VW���]�C�(���8P�^��Y�G4��:Cڌ�m�c�b˳ x#x?q�PP7��?�Cg�]����V�\��ᣲOQy,�`��.*ӛ����2~"zp��x�콆
��`�.܅�<˭.����#f���D��E,����"�O�E;���E����c�[��k>,�6��k��������O�uOj���!SD�)��FW֪�f�o�J��Ǝ��d��P�b��F	
�z
R,0�@M����&Yɛ�
�2"%C�Y#i��p��B�s��}���BK�l�$���B���u��5�E��.s�XJ�|�bϓգ_�n3�,Bv�4�Zd7�܇?|�/����\�@ӕ��[���h	�D.'��O^�N0�S`�j|m��1[Wsm�(�,Ij�;~��!?�>�<Q)����EM��ڋC�j�~��
	�O0��e�����T��� y �`���'��˘�˙�=�Pm��I3��ɬ�
g�˥�G�ጭOK�<����ǕX"�B_(�����P8�Ჸf$����ӊ����s���{.��Y���Є�����Q���X�S��4J;�>�������
�]ol�\��`C���`t���F0 0��t_��BeJ#E6I��:&D�.����IQ����6�L̘6�a��c����D�b�f<�~ FlƆ�O�����^V��z0+�{
~��EƠ����������Yt�-Fb������j�~��v7�c�,�g�ᦰD������/{y#������#};o_�b���*1�s�_��!��BP-���C)%W}���S�y6���(Q��y:ڎY4�]<ES!��H�	J�bhIY��`d}�Jo �WX� �U;98�ǱUj�z�%�ܓ"�Х���-�<:=��������H�vG�D�5O��߷�f��02�O�� ����N&00w�O�\������;~+TK�5�r0~!-ZC'ه��>���2#�K00W�l!
'��%�Z Q�l��t�I:�!�h�8Փ ����!��C<	��`j2`w@u����J,���h�.���gTk�.�&�I�q�3|��@���� �3�(OP B
������ꕯ#я WI���4�qӣ���z�X2�+R~��H���t3�n�h��"�#�;�>���*]��d�r�2]�N}�bF�) ��P��c�/���L�;�Zw����@R"�+�Xe����5�S0ǺB� �``�.N����_�gC�������,��#�0���ۤ�5M�Q!5���RN�T��$���2NRE��c[������'z��M�@����T��h�)�k�Cy� �:���:��?\t���;r
�6��mL��V������R�\��Ī�Ar�
���We`�U)q"������{>��Ȯ��d�HR�zI���7c���*Ǫ"���9��%����F#��9���86�ΡKr��j�m
�]}����B�"��u.���8\^����t��]b(���JT�!*��~�0��*���-���H7���뵔|�j�A��Qe6�"�(�9�a`p&�s�؁|5P{�N�3�!�!�����3�)E@���|s����B��W�;!y>u'����@���ZvQ�u���H4�Q�%Jߥ[�Bv�����*���e�| ����<�7���C@�����k/,�7?�I	+�\��'��2/գ#�oG�8����7փ\��2,�����mj�+�e�~���v�)����H�:G}mE���- @�vh��c�t�~��U<U�-��[g��]D=+.�d���_�g�4�C�6���$
�����>���V�ݤ�٨P�H�d��u����Y�͗���h�����<5K��u���6�ggF`�H����w`d�U� V6ź<�ǀ��5��cEH��K�,Tִ``;��vE�����
�ε~�Le5{�V��s=���\4WE��ǳ�/����J��b1zP2�]�4��*�i!{�$�T�F���ŗ��[�(�|x�OtC��ލ j���D2'㑒*��vc��{^���  v-*�-�㈌�^E�Pk`�=w�e�ĥ���)&��(��i>�|�$�3�.騒��w��� _[�&��b����	�X��2Ϭ&�*�ӵ����+R�=�u��
�'Y��ם�7互�f�kw�����os{�ՠ���*���1UB���]��������&L�!eX��3�ar�M-�,��e��A�o���+Yß���T��3W��w�'i�{3�i汗f3��H�����g8Qjӝ(���{���[�.R|�I�����}��B�o��.*~g8�w�^�r�<�W�Qb��<�d�n'5*ǿ5�����B�6|�H�PK�}2��8�����=�����Ur@�z�7\��Wɵ���Z9�ud[R�Yd�C�'�#�M����'��g�" �3�6�١J[��Dm��w}�t�dM��\��ah�!�B����o��P�����|��B��x���[�&��4���Mp��*f|K� ��b,��E �u��g^����[Sc�>~҇f�=hⰲ������T��� ��]T��H��!m�>����#��%�͟<��z�+��xl���Ƕ�\ P�a��Ȁlrq��b~���/���#�U�2�cP�x%�
��r�}����K,��.{g.t5ݿG�����59w� ��x(�X��f�N���bh�����U�������h+o��2�mWx��l�`�ėUD�ͬ{�C�@#����6��-�򏊑6�1|���b)����-�jk�����Kh� �u��U�5���vޔV���G1v�ّǐ�I&Y�>�h�遼V�4p/V�/C����XZ�r��#��ps����Z�qE�C}H#���݃3I�>dy�����y�Z�m������H#��P�pE*��ɯ��w|b�eW�ʑ404�������·���	�gĆ�Tg;�*�	D��n3D��@�,��4Ѷ��	݌iq(}�@-=9����m��w���X��a[���Ć����4�'³�W���g'��Cl�g��i�w`�~�����kd�8,& \ʰ��5�s@�l9o 1>hDF�B�A���1VFH�FD�8N�����l�'u����jxU�ͮB~@4O1/D�b&p����[���W2ubq;Oʵ(�ǻƢ	�@�A+���V��`탉>��P(Qw�?je�a�Q�e�MP}�9)�k{�n��YyVS 蝳Q>D��9���9>/��H�3�5�Xo퀌��vH�珟�����:a�(+�>�z>Ap�0�.��?�-*��0Ĺ#�!����S��+<M�^�z��MJeJh����]�wWL��g�m�} �����K��<�8�b�F�	i��+:��=`�B�8nP�Y���A�|�D���Z��D9��I��$�B^ӻ��`����E���	5�N7_�B���Ti<������~��Q4���Pk����/�����G6 _�5�����9�C��aJN-�dE� J��?����Jt_�Ӳ~���oq��w~U��>ԍ+���?�_��){�1*f��ؙ,.�=�Rx�K�>3!�\+��V��ZL#��*JH�v�bcU���l�Qp����i�X�N������X��*%��͟�Z�@3�05�-#IW�����X�},���2�6�:�Ĵ����������m�W<q���	?UV�K>7�#%��v�N&�[�oL���1I����A�����*p��g ��^�����$pp�ɂV+j�	����=pbL�5�SXq\��J`H���(�f����0D�{�}(���_��L+���נZ�6��y ���3�
8��r����y7 ���Ǯ��PeH�5���	���������v�6�%�$�����%iu�'�9 �8��7�ȯG�R�BE��Iح#?��o��m
��4���ph�zF�?�t{�oU���� �Ƥ��^��4wj���]֪Mz��Ƿ�L�H�>;���L��]N~�x���錘�L"ꐫ��IU��e�!��MrtG����������[O��tZp�L�ٻ��X�ܪ5� !Or5������lAR"�no��f.)��kĿ30����hQ��]�O�����yU�HsC���#���7�=t���~��.��~|y��6u��}S���|���/;Jy���j�=z�B��Y�A�f%�,�oN���.�K]~���Q_`?�4u��J�M���f�M�)c`h2���{:<W�W�O�a��=iT�h�c�u��o'�k;
��|���?�;�8�)�g̱i��E0�,I8�#�#�F��q���9g��<��8���[�$r��3�h���vd�������ꜞ��]����P��Ta_��̕���}����LVx;��C��>T�';��y��::lb9���H`2�,�]o�i�&�kk"�#(!y��E%,�H9;"�4bE!����(�2C�^$v����Cl���������5*$$���,�;�|;�uP�2�X�����@�'7�����rC��OA�-�j-�����R�m����7�/��6mW�-߉�״lW��v94�}�Y���T�:�����k�I��O�H!Ju��C�zo���uߠ �n���[����V����#๔Ҭ�η!4>�sD$�`������:| �"��_UK�[���{���|�7���7r~��$V�__����,GU*�%�����
�ABp�Q{�o�$�锦��Xd��`�j�[��9[`�2򌸸�ͮ$>��|s�������u�>I�̬*�O��ĿD�
�E=���d�LԨtcܥ�}�
8�(?uv��+K#-(�6��6�t��T~����M�UJ��v�۰x:@�_- ��)�L~sǧe�u�����V�	���$gv�C&�0Z!����� �
!H^"IL�l�7IXF"oK� B ݿ0w��b|�5ṉf��f�/����ad	�5���؟m:�}�R�k�|:x��oTlC;�h;�ku�6y<z�?��Cs�B��ՠ���׊-jq�E=�Uּ�̀���ֳ2����g�g��a_b5�I�@�fue�r&��%���Ⱥ.�<�w�q��bw�"�l�x���r4oǄ�#��O�I�i/���N��Y�OONsq�U�B��^�u���OE.��{�2Di��\��7�$ic��1��-�d��4�6����K�#�[V�'��~t��X��ROX*=��<���oP�����r�;��6zp(�T(LoQ8�O$�'����e��w�:��=%�>�f�>��F0����}۝nv�@�LL�X��{W[�BƩ��'����Z7$�L�=I���W�&Pߨ�d#*�����I7S[F��7>�E�-���A�D��D�i�SR�Tb>����l	�i%E��y��բ�qk�6�3�[@��n�LOSC���;����^-'�/ߤ��( >�Dn0��e���W��{��NWL�Z��3�j?�4�(?Jt�E�V�ay��=H��0� �*� j���o'��c;�]>�\�f4���;�n�1X�vw�;�~��G>ʔ.[�n� h����M�⟨�j� =t=t�aE��<���Ԥ�c�z	��];�Bʪ�S���)��&��H��U%��8�6��SL���Lظ�j��{�L�aK5����Ta������T���
M&��$>�^vfu�+�Q8�3ԶME:�L��S7�X���JNrF�4%f0�L���u˿!��-���-z�>3�
��/ ���BW�m�S�F���C�[�D��P%��L}�	=n�i��s�����;�*�L�̔^���^	�d�u%v�Г$��U�/��f���d�����WG��,��s�R@=��u)�oD�b�Q���(�S�)��[�]q .��'ܓ�����J)�H���h*�QE�����(sd����Ht�G`�,^3���K��g�nMy���z���K&��I��N:'��Й�F���w�W���C������O[w�;[��7�s
u��Ո��%������fђ�ʳ��c�O�lm�C�l���[l��2%�����AN�e>��h����q���;�6��E��(#�?���������6;�G��3��yyH����e���S���U@ز��d�e>�?��üR�M_S[,ӁK�-��{{W%an�
B�~��Ō�6���*%]�,Ԋi�S�Y#o�ĹQ�����mH��sId���lI�s|���ɲ(����sya�3��U"�X��f��.�:P pޢ��Z�9A���jV�X���a�����j>�p�f��j��L&�f ^ȟ'ᏚC�,����b����X@y¹�<�;��3=~��"3RX���!�ڳ�$Ѣ��Ü#j�W�~�����n=�E��5���^+�o|�Y������W)��(���.$�Q������u@m�V��s�\��������wO�ն���Vi��X�g�RC�|���r�4TE�<V4��L�zυ��x)��B5[ei�2�:ob�u<,	THL�r��^��V����N?�Z�Z�b�^�N�L�(�~�3f�5v�C������k��	P-�=b��PU��/�R��E[�	���OG�<���/ǈ�Mcx��b�-������Z=nbHvY�1��R�5�'���Ha�e?�n�]�Y���CHc��r���K3(Xk;K�:`F|��QA�7A����.�ղ<k��G���W̊8�0�ކ��D>\�>��^ց
K!h�~�5?�:�a��~��`��8���Y��^�?�0��Md�c\��JI%H=�_x� �@�@X�����{��E]֝�>��z���9
�>L����T�R�`���K�y�z�*,�PO�x^;����ݫ E�O]"�x�K��KeE�c��D<J��`qz��ݰb��0��lɽ,��O�q�KQ@�w,ec!w`ǩWҮ]�i�Z5L������,� ȭ�Q�Z�U0���k_�~9��\WI�!���͙X�>R��!̝9��AXW��Ě0�W�-���4���& 1tr��qJ�q+�f� 7LʭbS�Ǻ��@gz�����T���Fq�+�kI���u)m�2WgAt��l�'*̼��p0�+Ѡ!t#�������[_��IQ�1xu��.*e�؁�#4���N�f.	�3���z�^��'��[�vV���l�hg�}a�3�8M���;�O��!�g|A��4ϔ�:Z��B��*��\A�U �H��a �X�l7��iu�F����UG��o�2��Jw��(���hj�_tBt0�&��ģ�����ڎD���e��>̿�o�X��������K�ǻ�F^�?�8���m���:Fe qUQk��2>����ˬ� �ݷ#�����Ho7[]�m5r;y���<��VFe&��c�hŘ'�6��~~b�G�HM���;�����9Ng�q�Zj�5��<k�I�
�=�yPy��N��'e7u0Z~L�Bv`��B��w3�f�	��/l1���F*�I
!M/\c6�E����q�$Xy#Ӧ�Byd��dQ��aZNp�������=:
$(�����������G�Z�v���J�"��oX`,c#2�����4D��7�V�p������OF!������|��Z��b[����v���H�he �*����	(���Rm�����g�g�����ǅCe v��9�+�iK�B��m�SNqF.S�,RJ�m���	���Ƀ���!���N����{?���"����ڣ��E��z�J�t����1��D�!�2A�#Bt�ob�筺��1���/C���-���/0�,L�r5s-���$����n+7��J���r�Y>m���T�jbm�/�s("
WQ�����ĳl����pE���i� y�H|az;���6��@B�A����'���}F���7�x�J��-���j��n�������V�����+GnZx��6�'dX��?de�$v�9��G�v�C������36$���_�u�L�����-�%��ğ:�a���ءwJͻ���ａ;0x�a��8�՚۠n���
q0����d�j���20vdl�q�g
Zip�G�����>��F�&LF�N` �pN]_C��� K\ۛ�c����I���>���$�Y�8�7j�;a����AE`����2���_6��S�W�W"D��>j�}z�pS��{D�c����OJ\mL��j2:b��n��©��C>g��裡�
+��k�8�ր��S]ȻdO�aYl�J��od���[D��VY�ˮ���o>^l�%�*'� �Wj��ή9�8�o��1��p�Y����hA>�l��>Mщ��)�KJ��>�:��z�.���775��v-�������l�0�ˇU�,�Ll"l�r�S{�X�sE0go�l�v��y���Dr |N�1��Q��"�W,��WJA7Y����L��hlF�6C��fA��ZѴ
/A�z�<1d�g��Q�jMG�Q�0���x���h�k�T��:�����ӌu��I���r�l�3>�s���q�~���X�c�����ɚ[g�4r�B�8�{�vj��6]#��p8߿�?uvP�� �OV�O�ö�e��< �A%��s
H��df����^)_Xf�t~���%����TwͪT|�>{1��4�$�W�����}m$AĠ@ްP��b�1��.�. ��j�XNAk��ѳb�et:Z�i_ՐF〱��%z<�=":��O��t��
���"P����KUe}e�?�j�,����Ӟ3و��_�lx�s���dI��	8^h����7k]J�Tr�b9����']�<3�����}&x���5TsUa�����\Q�oa���b�v��;,�,}�%�
=��R���d�e� R�犿1�A�V��z�\�x��S`�(�O�ജC����6���M����z�xK��=�?6�U�Xm�
RF�wh���%J��S�A�م��e����+K;`��HJ�)1����2�)�nj��H�����0�v[�wm�x2��d�;t`x�ALv���x���
L?QI�g�ހ��d�'��f�Imu[M]i��k�H�m9Nn:H�5 ?�mܔ@H�vi!�.���1�T��|��"?�*][y�U�[��3���5E��` ��h��Q��s�j�Ӥ+F�kb����|έ������cT����й��VT0 /�t$�9��\1���N��q��hv��LN����$�0.�C���
��J��e�����=}�>mx��5��_�^�h
ӱ�%�^�ϟ�@����`�a_����o2;�FBNT�"�d���t�a�Wꪪ5qVC�_���?9��� ���:T��i�Ǆ0[�~���.�D�<�X-[&KZ�J{��~~�+C^�[�����#$Ñ8k���A���qa�K"�zk���޺��E�҈���~�׉4i��f�%�ݑ,�cgs�&���	�^�v)�HU�����5cZJF]9���3��zN�������ΐ����y:	K��v��o<��>Z�X�t5h�mCʡ��������,���eɾD ��)�,ҧ�8ڪN�'�����9�k��F$�7
3M(Z���a&�꡼5�.ݵ�C�����De��(&݈;���ZB@T�Y�����5�똟��i�i��++�Qin����#E:V�mD�p�=����:�?4�6�;��p�E;'}��$�<줅V�����?����d`;�~������Y� ����ك�W�b��{�i�/�z�V�\,�{0��Y�*Ri�<1`(��$,���1�3B����R��t�h��,�u����E�����HD,9Q���;�t���%�q����) ����~�0����߁2�<˓.-�me(�Iw*5SfM��b��a�u`�/텴)��Dzd�Z�F��~����\�óuJ��e�c�u����/�;�����V�a��&0޶[��ps��Z3c�[�.8�e��{�I�mkm/��(�»�WY�Uvx3�4�Z�^��r��������}N��)ٷhzM���XI9y�C��5��F���x��⬏�wkC=��$<قn������c9#)��5��?�򈭦�df��� �c�'��Ro�Lʽx�ּ��c){V����7���;|�_20��c�����m�a�P����#{kRF\jά�nG�E�"�N�u��C)*�s���S�ʄ8WMl��j�T���R����i�d�<��z~���L��"Ȱ�'=��Т��m)�O�\��}OVPgD	Y�>��93��'ӌ~
	��>Xb�h�!���F*E���-ˋ�^Sq�`��Ѷ�t�&����5�|�[4�$�Kb�`u� �i?څ���e���'��4���Ӄ� �î�ֆOc�ݠ� ֈ7e��`����vs?/��&�9L�WS�˥C� O6
��9�+B�9v��@Q�G�����'���� S�����ZF�=_��U��}x�k���j�L�)�-���T��?��g�:��-��i��ْT[c�
����!���}��Ϧ����;�̊�R�5���m�̕Qa(�KWz�2��Z�\�n|)0^�j���Ce��]Meج�.Sn���[�Rk���[�.�X��&�㘱��S�[��垼�.����x���ͯ�1�� ىu��P��==�5 ��1GG��0׼� ����,���aB{�f�";��}>]�Vl=4NB��էU�� d��x�|�+���L���%4wJ�x�6/��n�R1�m.S^z5��-����m�r��t�\�d  `��7����VMR�%���C9�>?6lK)k[�N7��ؘ �?�p�m(��ǁp�Ռp��M�S���)��9�*�Z�1ٓ��2�0�#އu%U&�c���$s{%u�B!�u�t��?x�='�k~�O���!{��[�[ '%�9�i�j!=��N4���g�>�)YD��&�EϺ��{y�a�d��?Y�4�U�����\Uh#�V�Af>5��3��Jg�^m�U�B��/0H��H���_��I��WYp)Tw�+���d5ܚK��������2��k|'�s_�f��9d6�}���*����[{C��;�y��D�Z��!����)�q��<�/&�x\� �2�
��6$�i!V�6?�� ػږ����sH(	�a����3Z� �f^lf�.E~���ii��O�� 	7�V��� #�3�Q=��"}�,Y�OXb�H�鸽�вӬ��ԙ���[9b~�;-�E9�U�� &+ό�t������@X���h�1�`��I>7�e���u%铜p<f���jf��6/�?B�A��s�]G�[m@e�A)pF��]�bJ2��J 6�q���%y��>=�|e���&3��F�B4�!����,�GK�)N���v��Q� 4��e�,֎�х��u*+%;�ٮ0�3e���".k�kR"�N�*-�XQ����-�&�H��(`;�:�n�
�eՒ���?ɍt�B� ���9T·C�MB}#�S�0}�]\Q�Q����B������ Ga�X�&ϩ��΁�Ga�J��ᙗ��r�P/2m�J��X�E�+d %�f�:��Ro6�bӼ�}vN�&�EU53��b��Im������f-��%�j�ԉ��<s-�S⛒�K%W׼@�+w�/c:IO3V�)A������ge<�@]�MY���%I?^l{�`%������z��!c6��c�5/>bz.����,|��4���x���e��а"�ӣ:ʖI�Q�E��6:51��5gk��o�I�rs������F|Z
�T(�����
oU�E��6�GO�jZ�@�q���zY%)	�ۢ�[<�|��L�L����9̗֯��n�L��mL�����)��������bZA��njܶ��T50���i�D�����⛄R��39�:��g7�z�{5�y��(�<QU��ɓh��������8��L��z��m�`D"/Bu@XE������@rt�Zp$���'�������:^�����1��� H6����J�u�7�yp�K��6"���!U��9^a[V������%~��|�ݟpk��JިIs)jk`o&:���Em�G��,j}�
�	���wE���-����e�p��&�v9%�.����yͲ�f���������/��7`�~��ꚓ�^|;��A���G���\�e������쓎��Aʴk��VV�Y�e5W��1=?<�w��4_3��@�+���`F��OV��]���6�F��NYߐ�L���}����>�K�����w5-��T$�:�/"{�L�w���o��QX#��Ў�A�Q���[�"ϖ�y��Rd$�_^��^�3�~�孈��cl�Fk�9��t�V�(�(�"�*�x��Q��K������3-y�e� }��`�Z���P���-T1�,U�ܽyM�M��O�@
�=��U��(nP��D�P�/[E���S�Ӹ�jz���[�o󱇺u�!b��k��9I��'���~�Z����Ie�#ڡRn�P�qiY�HoS�ۡ�ꚠ�J{���t�w=V��d^���m}x���8�x��������������.�7�܁���c��^	|A�*���<n|��gz��Uz�_l�m�� �I4�ɍmI�Q�H�҈��9q��hP�s��h
E�4����Pd_G�J�׫P��!Ц\T�0���w�}kA<�����O@���|AƢm����u������6��}m���8��~^�I�z6`}����θ���@���vY�a3R�i�T�I��2.��C�^ ���iF�k7��z ��vʧ�ԝߎz
tb��FCc��rϖ�Y��,�9@���U��0s�m���GD���%4���y'$h��RCBr��3+��7%I��\�EA"o�l��@��8�j#�q�|ۣE�R�	i��N�h~�R[K#(����"��i(OW�A�-s�7gQ�0��"��G�� �7%ڡr1H{/:�z��@ql�}�r�N���\�v�@���P-mFE<�G��U����Ͼ^��P�qy�-w� RK���`a���j��lH �|��+��Њs���߯~�1IљH��-��e�k� {��o�����r��\�/�u��=\�z�g�ԕ�� ���|�>��!)Wu2���#2rLZ�o=C����j��Ǡ�Ħ@�.!��m@^����Y����AnB�ͭ�(����3?Y�5${��.������b��$#,=��q氢_
��0u�DBM���3�i���/��-%r%�s��1�������%z�T��Ί)�[J��
D{���!�.��.� }3�-/�e[T����Kk����)�|��G��	���PG�Ȁ@���A�8� Tph6��&������'0t�D�)�ך�+��}u߼���ٹn���9�
�Ux��W˥|�F�H�p��vC9����Bx7����Z���B�)�LH��/n1�7uо�a�c����~��7xp�]�1�y��g!��*D:o-�g�f���!�	iA�f�AZ��ў�߾�&�S|��!q84��`µ4�l�M��=:!�~e�������L��R��f)��PE�v�Y�'w��x;�G7��$*��X���p�D����K�S-���QH�b��0��Y�wrz��YS���9ӡ�h�2�*�H{�41f�{A��8�r�~+��LK?��e]�`Y]�P���'���7���C�%�ˑbT��M_h�Ћ� �)�}�9��f5��U����7�87=TrI5خ:J���;ޙЭ�H놢�Z�%��2�7O�8�%�MPv;p-$�j��LYVJij�����z�R݄�8R�GF��T}�n$@�J��F�z��%�����~oU8#�R�^n:7����W��)��ƹZ�'e���5X���E��A������_�̠)#���d)e)ݶ�	,�P4�A(�j\,�4�^���ޛ�W2:��0�^Ԟ51Y�ƈ|{u62�5_������U;[Ja
�*�_�V>�}0��)a��1<
+��{�<A.*���-�3����<:�ͧ={�Si�e�T#�S��!�i�q*�<��Yn�8�QN��Ĩ�`�.\��	�hh�0_���'`�)W6W�à/����@��&lUV�{Ŗi!ߑ�I&͈�;<�Ve�$XxKXgM��.�"��E��X�V:�elG��H�$�h�7!E�t��v»��z����ˊ-J�ْ���|`��f��DWX	�a�y\x���uO�;y�o��|�_F��*_�Qn����Ëx�<م�2���ւ���l(��}W�+�'�)&�!Ա�4�pl	�4�B�W� ,@�5�E5Z3�B�r�	+ ���C��$uA��QJH��Q�W�f��/Z�W���2�f����öP�lr'����:�]m���
�f�n�l�[����j�u]�F��r��㒑���<k{��f���o �����-�~�'"�͸�������2�����q-�YLS\)���6��,, ]o�����Z�IkX�+�R���J��8g�P?XC��+�Ց�םa������h�aG\�-���ނ[��2�[��iz��T�?q�r�c|��^mۇ}���vށ�9+S���#Z�+���Q�C}��vV�$�4�$���T���
�@}�������?!��*�Ci&�Fw$��Aq5���\V_y��ҩ���k�"�'�m��#څ	ע����R>D�^�6��y��(�W�Ff���+U;/�f�9ZH�I�r4�����E�����%��� �%���6Q����{M�gwXee`��S PKޟ��P�S�Z��ɬˮA�+���
�+�A�o����e�����R<�s	�lɏh��`���ή�0c�%���t�Y�̫d��*��5 ���֔��Y)2m��	���Dz<(�ySq�a���VU@׆�_*iϳV;$�e��s_�P}DbF6�vJ�W��4��C��[^��OG  P�d�V4�s��F����x�K�djg� >��8����x/��5�͊��Z�P  ß`����`u_R�]�*�_⑒�{�V'�#g�x���+YXa�i�m%�j�d���3�F=,^1f��K4�����G̖k �N���x��!�6d�t3\���ۊ�(1�F���T�����*^��RP������>��U\�}9�'�iK��5�(���@��.��c,_�w���o@}F��n4w���e�������}�I� K�cp���:���;�EU;���Q�0U�_DU�tRzJ�y�(���)�}��-p��qݴ�.���Ŗ:
��Tx��t�S�w�'�e�(����Ӹ���7{}$�

5:?U��;���]vj���6KV���SZ��v����2sq'�h���Z�����^����k�kM����O4�/��	���dK���简�����ZE0�Ҭd��f�}B#� �C ��3�	�GKoY�$7I~�����a�K�(=��@*�g��2�}x�o�m�g�L��+����p}Ns5Y]]��y�þ�6�7��&i5�5�	��l��:�$oK�,w�{.������뻴�_�*wa�j�ٵL�3�r�0ucR�M����̋���Y���Ғb�;�K蔬�#���V��L��0A��C�E��Z�ь6�X�R�N��SG�𖚠6'��M�R��vJX�v^#f_���[u$���UC�Q�㢽 �0�@A��'/�bVX�����k�)Q�ɂv�[V�T��O0�"��3�cݐĘ������9B���|�^㻷O7�Z�Dj[<cyc\|����M�J���>O0^[Аӛd�"څ�kᕑRC#���[��W���4|m�0�	���2�İ�ژ��:�5� ꔂ��'�V�}�"m	:�zi������̤��FA�/�b0
���O�Nd-�N'�BF|�d�#���VKn!�_�+�L�{�`ZA~6�3�O	�6�E}	�P���>g=G`���S�C�6g$�d$�im�����+���\GV���v���Ho���"B���mLHt(yԦ��cc����n;LD{�MW|%䮪�,7�^�hԽ��C�F�6����[�Ţ������O.�ç(f��ީ� w�稵�|~xơ��ċp��w����S��
�Ɩ��� 3�'��>�Z1����RS��X|��_@�~��ʴ!����k�8sh{�o��`V�L�E��;S�dx]�d��D�`_"[�Ѓou�\E/��q
?G�y�mQ����,�3�"J@µڒ�/؊��_�^��7"�#�?�v�+����@�V��T�͘l�!0p�F�m�����	� ��E�W�<.@�*��']�����h(�n)�]>}��r9�#�g���RZPg�Ƞ˟�i�]���+#g�T[�}�&���'�V9v�xFH���%��k*�&�63$`T����TO��,GG�P&p9��]�z��S�ل.�0L �A��Ѯ�Kdk�L�`b��>ֹ�MY���Fw�>kAN<��V�Ħ�ON5��%J1��{iC��`}JU()�bB�]"GIE_��m���I�����{|�x�gSu *�g��U����i�>�3�w�ID�D��7M_Adj�!�wE-�w����,8��U�C�!�ה!4O@�Oiu��ۂë���O���֏��x�5� �ʗ�~�[}^�]J�� �{���0��-�_�͸�Ӏ�,-�1@D�v�gW_�F̀�_Z�̿�^]��	�I����.�S�]�-5DZ����=�EïxPF隚��ˉ�x?����a/���$^K�%�9�@8�^W�D敉Ayn}핾���z���9�ԡI}]%�e~�:���<���~"�ʨ�1g������΂�0�ҷ<���P*�]j��Ɨ ��KRk�*1�) Zo|�q���^��V/<k8�pq[�h�{��%����Q���%� �T{�-cj�ЈY�&�3@*/�j�C6X%��onr��O��,6Y�pi��a9���{b~J[V�PCq i-R���o�T=��V�ɩ�2�D ��<K�����<ǈ��r���υ��H��F����A��T�v62��<u���Pge��+�f�S\�+ag�y9�X?sQƻX��"��Φ��>�$���
T� �M�o�l���N�½�Q��|e>�%5i�����ա���ُ��]ہĘ(��B��p�i;/Հ���qU�2�~�WF�#�C¸df�ŭ������8qE慭�Ԃ�����V�� .||��Z�Ձ��M���ޠ���)Ԉ݊�M)��ٚ�KO����>�v�>���]�T�4�p�}�3�o/Ѓ۫2q��Y�W�nmha_��<�s��q]�;��#��3e�07p`�L�'n��R�!�D�"�f��FIb�b�N�ݓN��!MZw��
��K��]wvuv�H:�y4ڢ�bbA\��LЭ񙜸͈*lpcڋ1�x�8��`��,N@����Hw6U2���ŵ��s>4���� ��%��M/��X���-�F͖LG11���\6����}z}���zwi���'�W����Ʌ�A�czCҚ`6Ê�%�3R7�_3����(�}>����:��Q0I�z-FeF_��랴���6S�	��}��E�t4;2���ąN<9�)W�Itd;�*�J����M�Ou'6R
#�r�n�&�(���a��ZjgJ��'�2eh򅓃wM-��|],��Q�QH���\T���f���a�_���"��&��G�֏BtG�'F񄦳??�W��dc�>��1L�L���w�O�p��72y]]�a<e�#]G�a��!rŃ��H�����eǝ}�)�������D��c�A�.!�]��2*� ��%�p�K�pj���H�	�js�ߞ�S����'|i
M)˧on|r(�����Y�rC�r=x,�{��!�p���0o8�	P=Y��Э�O����1�_�����M�l���������$ƺh��[����1�2䢽p%Z�~Ɂ2�N�8(�OϾ�Rî�'Ҭ7�F~��O�x!��Ꝭ����;	 7�b&O}��"�{t+$�rIt#U��(ů���vZ����� ݹ��(�r�Ƣ����p*<�D�4š(J��!$>�GO�����e�����@Q�@���xu&������NI�u*��A��&�;O�LET�m���"Np�.,��Z_Aw�$�s3�­i6�NT���͌x�$-g��Nh�y�R�(�!�#�m�����_M�ޑJ{�:��ׇ�iHP���?��}���d6��8�; �x����&J�T����Qߖ���
0g���T�/�����KS�
���=��3��ܦ����p@R���m(  ��w����l�k�͢��o� �UF��mm8�[���P�l�r� �x�#����N���0���2���`B���)E��D��LE�ǩ��>�@�����ܝ�>�b%���A����_W �nԧ�qd2lʝؤc��D
�P6���`��,6����ːC�m9-t^#.��:��>�n�-�!A",���~2$�3,"�uK�nQ���Mb�CC=!H��L(0���}@谡�a������N�f�K�}/�r��I��B��M������mqo�Yā�(�����۹�Y�~���|��c���YS�?��0!�1����K��]1G��]M��Y���O`�[�]�Ky�I�7�Q�K�g����U�7�vN�qⳘ�XP���p�m��9�R�*���J�	Y~=%ҵ!��HR���a�˕nZ��F�v�d�
�L�wR@wČbGl�S�E�{R��N���'R��t�����8��u�wƯ����"á�Kk���I��Ti�k����xW�<ڥß;W� ��b��\�G�s�@oʣU��%��d����:ky�̆�(0b����jCv¢b�� �S���������Q.�-D�ּ(���IքV���ħv<�Lйj<"�g��� �8<��\*�� G�7{|�����������e�݊�ߺ�9E���������~�o!c0P&Lf�Y
$�"�߿n�fVw�Mʯ��0���M^�0��Q��sf?�GF5R�a>� ���,?_s��K��t�6�����-On��Qn{���U/K!��L�:�\��2��$���"X���#�a��Z�xI������ߌ32-��9V*V�ߩ�A��I����092��X.��>���Y�m�>��5�:@Pfi#��?�kb�/�n:�2��)9L�K��+���[i��NS�B1!���[��E!���]�V�߀�����\8sI�z����#/�N�U�-Y_	`��ms��3	����o�!/6O�䞸x(|����K�>��#<sW�B�i����>x�
*�"�)pM�mv!G�:�ՃG��~��ϹI6�W����L?���fu�G�!��'k)��a��ߡ��t�`�d͇�>�I�E_-����s���l�sS� 4��8�+��J6���h�L��I��xEW��2#Gz&~��A�j�K}$��~a�����鋍��6ͭib���@T%pLD�$����$)�lHHş�Cq��D[�\z=_w@3=9�p�޸.��{U������}�����H���G�0-Ȕ�)xNc�%���A�:&�I7�������Uq*3�PŠ9�P�;t-܋Ħ2�V	������׀&���szeF�P����F~�RU�V4�nO��u����ց��
A7n�܃�m��IčHP+���"U�f"�����3�$(֓I$�SQ�:f�J�̓%m�I���	D4-�h��kM�����GP�x?��9�����yuw$��7(���'!l�N�;7��ca�ňtd(�F�!x-W���Z]2o�M�g@4�ߓ�&��P���*}��O���L�/W��j1�e�&�Gt�:���CϢp�L7���:;��Pg�[ӊ����q�Pgs}�ŀ[e�������eH��S�,Vޘ���[�UR�e~f�
o���>�]����6!��"Cmh��Wė��	��M�*�1�XYI�96�0��%�,U>��m<��̹��������}ﵶ��XlN��+8���#V�$'�<6pa���T��Nz�'��ňpU.�֮���W�p�y��O���j���_fn�s�
���]�Z��Q;�ߗ|�0+d)3Mʹs��K�m<DC���kOB(Sk�U!Z�i^�L��M7d-���|-<ϖE&���z}��o�X5�M��ˬ�{2L�"�噅k3�hه'9$�X0�iJ��@�37�R��ЍJ�]��XR|�+t#��R����e�����1�@f��|b�w�8(�4z�ѓ��_EK��v`�!�����{䖼�	�'~T[1,z}��B�y>��������e�끱��G��[5�|↴��L�W�k����&���K1�'�O���uW�j0�C�;��m��y��m	�*Nu�
d|�6�|*�!�s[�8�f/�P)hJ"�-(cK�2g��X? �s�[����R��[���O|.�4����Rc��˵C��k�$�/S�I�p����F�m!��2E��!��b���|�����{ؿ��E���"�L�0.���y+	��[����v��`
�eH�_na�G��Cv+�7Q��2�,�m�Cd�Y^F�떓ևG^�39ys�Ȋ�^�;@��WSKN���#3I���d�u`����H���5���({#X�~������Yc�.g-�� j�w��E��'��.�����Rx���c*�����N���k\�餃�v�"Θ���D�t|Ǫ}��w�Ʌ� �
^����;C�R�@���1#,�ɥ���&r�,�3��"�n��է�> [r�=�;4����M�����c�&���g���&��S�N��V������q���j�ˏ���%���Q����6d�r�����[��I�������g2mC���t�������<NyA�ǺY^6tש��*�Y�<Ԛ�̎H�:�L��UfBo	��K�i��z|W��Y�R�{⺅Z�+�H�Q,&���fP94@��lC���32e ��	T�tf�KjeW#�\��9�*�<i�X�C��ztC��|�z fx�%�Զu7YwW�Jbc��kf[���=jJ5��	̨Y�PPOm��0����\��;%��a���8a����kr}�=z���9}$#}d�M{�l��NTH�A��W�����E�Q���n&�z+]��!l�Gݓf��^UƛO+�bt}ޙ	|��U�z����&9>JvE�� a	�EB"�v2&���{k���]3���i�.��{@�2,\�s!�UA�Y�n0l�Pb��w-Y1�1��Ҿ��O�
��3=�^�YKՒ�wL�����U�.f����G�Hs?+�M
�� �\j�k^eę�E|<� B���ZE�Kf�$24��OɽD���诟t*QơEA},���Z��N$+rܵ�v�j��!.�C�C�d���P཮���S�B�..�� ��=�����c'R�&� h�3���z��8kj��hv$3Ӱ�
�����N_���`�R�q\��)ث�JN�1z�~��?fZ��YH����X��Ju_�ݞ迥�4�)���n��>Ad��<�6�� V������:L�x�=L�=r�ߦ�� }r�&8���i��V�$��� )ܥ�s���u�֧u{�E�_��Jx�@����� ������5����R�O�g���Z[�P��o���E�$޽
�0���l�_���C(����������W��,+��	��Ov��șDә62
\7�[ �A��A\Q��"�K����<:��ĠrQ7�v�� ��c)q�Z0����o%�=����ِۦ*�3%�[b��E剤�F��C�B֎Q����~ 4�W�{����P����a*��7U��[���ſ��ӑ܄�P<�ʢL�_����>��<�!�G\�?�����:��eW%/.M�Y醖6 ���<N�K�$v��F|i0�vȨ���o����9k�"[���L~N��y����E��
�x�OC"��OV��3���}t���)�m�fIi�k�����J��\L�B7������������)*�}8\���Qv�����QU��;Ocns$-rd�t���܊Fq�����47\ž�F3ȳ����-����A�M�n���X��?¸��f�љ�DB�@:��_�"1���"&Gݗ�{Mq�V5�᥃�_T[�ti/~�ߤ?���!�1M�bH���T*�R�,��BT�lbt{e>柞�o�*{
E��.IN-�D���sK�7!��'�4�|CWY�"32B/'ICz���[���Y/��xv�&�*Nڥ0��E���q*�#�ǅ>�w�f$��n-s�f��l�#_����/�Dx喉vS�K�L��ϕ/�M���0��/h@tzD15��{��Y�%�u��g�3���ǆ�D�����}���0����z���/�p韎[�|2)����5.�����Z��G� 62�r��z,!�$6��|��s\ن~��n  �K�H��:�&����]�=�I$�jΙ����9k����P�������^'��0��љ݀��(uT���(�ؿ�����d��@�b�h8R����ĀS���ʓ��ԑ;8�K�>a�AL}Ż�3���4���O6�s.�tF�؀��4E���J�*U�v@�P���ۑ�lu퍆��H�phLNy�6�I�^|���-|�ċ�!�#+:��i�w��թ�/$z��%Ċ~b���,���q>��IOH@�����r�M�L��.4���� �h�����+z�j�U���Sh+��Cvb��w(��)<Cd&V9A`�WL�2��u��D?t���@_�J��?
T�'�D2��"^@��l�rDUX�?	ϙ��x(������Ū�:�[��Fh���3FA�|���｛� nȳz�7����!:'�v���J����=�����껙Vsqo�u�,��炭����՞�|�+ٹYX&Z��v��~48��	f��B�O�Q���=h;)�����H�"֘���߻�ϥJzڠ,�y����� �k�.���8{�G� ,|�`��,�yg��i9��(ʾ�<�K�Pq&���Ϊ�Rz���&L(:T�{zΚ�����%n;m<c��rB�J�p������q���6���(��0U"Y�!
)�Ipޱwj?��P��zZ
f�}c�Ùg�YrNNI����0�_ĀGY_!h2H�%J��n;9�w��Q����8�aV ����%Id-������	�}nN9�o�3[�"x=t����
$�蕧;�?�ۋ���f}_��
|r��s-=p�񝛄���\�O�<�`)f��Po|Ƒe�1�X^�?�@�(pr�Zw����Տ�-+��8�9d 70D4.��u�\=���}	~|c3�Ѐ���F�ۆy����$:)��`��pȶ���h�|v�{��Tԋ��P�n	5�����C:��?�ἔ�*}=�0<� ���1���#VX�����/�e�o�Nj�e�T�E6t,f����	��ܡո�:�2���>�G,m�	B�\ߛT����[�ܰ�X��j�pµ�n����B��N&Ho��"��N�8ǿ�-��2�yb@b��"toӢM,A��Z�^ᜯ��b��_���}l��$�#�$b��[m&�I(��h1b2���׾ٮ�mdġ��8f�~��9������(Pk���X�=��*�����^߽F����&m�4�&�j��-!���l��ٯ�2�Ɉ��/��/,���Ҟd+RNj}��Ov�2��ʈ�l��}�f���؎��w����b� ��8K�Ӡ�O�F�� �0�I�����#;��ƶ�
�s������4 -o9'�&mr����k�ڣ� �{�e�x� ����0W���z��Q�Ւ����12��՝����>��}4�(A|US6��l��K"���vr��������ɧ�GXÖ-h�#�z.�ٙ�ZW6ڽ"OB#��g[L�OX�{e$޸��_���I
&e�����]�=mO�ŘU�� �W��9���p1��:�Ʌ�<9I�7�c~)�� �[P�i���$�s����5]�c,��q��V*5�{@p���uQ,?��S$8m�֋nN>[�T4��O������_27�JY?��A��*�{�̬�0A�����d�k�(��#�aB�!� Ci�Hס��4�L��i��$�@Lz��� x׏� ᄇ/�Y�D�C�]�(���F<�M��'B��G�,�y���rv�{5u~{q��Iu������%��&��Mj�9���J���6����}ː�J���n;Z���f��ᵀL�٠�� �CG���7���%�����KX,~U��HT�܈{�����u{-r`�`��W��~�@`�ભ�8m��	B�c<J5���;�93�Y)�m*V�~ %=�k�6��������<$M�,䫩�j����%C:��Ә������e�$U�#b��iP���z�$�9z��sR�K0��EĶ­q���li*���T`Cl(b�Aix����\k{I�B���r�%߰��{I�W���Z��)Ԭ�Rc@T0e�AB��wFa������}�����>���;�E�Ս,!���ԻBH� �X5+�p�w?u���ۜl3�bV����;�Qj(�q206�@����1�%�f�{�\g.w��S��]���>���rNV�|���%��0-� /��;��i7\��<� �*X�J�2I�p�s�DU ~V�������!S�#��dL��t���x$��L4�lT�4��S�QR2� P��Ή�Ǧ��{�Z�+>��&YW?�b�hm�r�U�d�PK ����`<�S�����!�W�|�0�&V�ٙ�6��Y����첶�9̏�ɜw��ͪd����E,�6o;��a�����~j��V��7�H��wv��ḩ6Wd�Y�I�m�:�q��τ�$GLđ�O��`dF��*����x��F�o^���'qپ��8S�fA�N>8-R�8p��H�JT>�6��2��L�益��	��:i�*�%ݚEB�Nm(e�x��G��+�º�g-�|�aե���b�K�Q`���J�9��K��K��ڷ$��)�Vt�@����H�K�F�b�"���b�;�51_����UN��GiY���wO���ؽ]���뻻Z�Ê�
�=�3��G���B~���uC�cu⍘y�%_�WO�~�����ݦϹ�Lw꒎{5~����CG]�c��#��-���a�~�~ጡ&�A����p�<��xdu���5Z�|�f��Z�/�%�ESbd1Ի5\�	����]�V
?��sEp�g����׀�4�;ޛ�Nv5A��?�X�Yr�:[�
0�*D{X�r���7�#�5��rr 9o��\#�'S+w�)1�is�;��K�ś�����]�-�Ҋ�3#Z���0P�����;��Ƃk��3Թ-��4e.�;�Z k���k#D�!,\�@�M�k���Lq�M���k��b�4�T���5�E]'�֗��>�:�����ů!DJr}��U����&rk��V?q@�}��dn�U�,�kzp�s�F�p�nF������>^Z-���=�H�ƺ**b���x��Z�mqd��жo��I; x����B��V��g�Ƌ*17���.tnwu�1/76�H��oU~�З��5�6�7f~�%�b�Z*�jq�0�;zȗ��0�e��7%m��,�w�\+�(M0Qf�@�n���Ux�3fIO��� $��E,��%cO����&�
뎮,3���,v�B�`<&�� ѯ"v22�Z]y��+�"H���&pU��rA xp�Ռ7���V�+�]�h{��"=9�X���U�|Z����R�p�Z#|C,�{VC"���~�`�Q b3ʸe���i�"�U���D�ҧsS��xQ�)���!5�Ep]
�S��x��u4J�nJ?f;~��16�R��9Ddc�����4��*[�� � ~s�\�lH����*����d�^{+U⮛�sx���J�Mͷ��b��Jڕ[Ǫ�mM�fU8��l)��:\�|�hP*�.��}&O���0�!�<���.X�S���4�0�ǣ�G"�9�TM�U���q4nj����5�Jњ��!m
���]}. �&�����n����&S�7H'���>4��H���~@bu�6�w+t*�QVrl��}�s� s���Y��spIm��4��?���<8�4,��w�+F�t�G�3����I����� �eP��p�y/�]�2��$��݌��y�Թ�)oۂx��N&T���i��j�������6(��C�w��m7���(�rԌ�~J�λ�ƶ۝P�gu2ܫ
��&r[����s�Bx~q'uH�+ߠ��CK;�/�-+�c6���B�K������{��8h���"����_o1c���_���aXw��%�L!U��2������P�!�u�t���2:�~\��ɉS�K�e��IPB��;���y52�$�x3Pu$XV
S_��\6�C�{��a#���5���HX��2���g������?4X�����G��C��KG@-�(���_ �	�m��ɒQNRwŜG��Ǎ#�|�L3jːLO*ݳ�P]`BT)5`1r��!��s�ib ���o#- ��Nm�K�a�����M�!�@}p<���l�RI�Ț?�d�g����Ge��xhs�_�ɰ��T�^���'�A�PPy�	wm�^��{9�I���`�쳒�|�Q��x���}H��&�[���=ߚ���Z�؛cJ���_Z0\�B����A�Om���-�,
�H�i��Geo�q���n��'y��H����8���}w�lb�x\ K�f=���*��-�2�$S��Uw���m�r �	�^�¼M���L\<\�md�v�8+L �aKs��̇�%��J�LE�BM���!p�&c��%m%�%���X)`PtH�]�ا��:�} (�]0�=IP@d�]�"�E���f�9,V�o3�����!_[ɿ�_^�aK�Um(��Bh�R[��O�2d�}H���%υ��]���܀]X:��=��-���ڈn�nR�V���n���O��r��*�����Mݣ�����3�:M9�2�M�@Y`7W�R5vZjL��L�]Ȁp�����LP������G�j=��w�PR�� ͋��ڔ.}�d���'�+�:R>94��mc���Z�G�;�43����Z��L�	 GF�u��ώ���!�U�(�'���އ�O��Z�c��š���q�9p�ɞ�εѼ���.�]���S_nj-x����D54��F~n������e�!wl=NH�5�l�
�9�7o��������pP�6�I/�B²k�N�>ԾJ~M`�~5��w�q�U2ĦB-���ѵL���D��O���]���F���v%w[o���P�q���o�ԉ��y�eV�f����ŒZ�,�Nq����o!����~Awr�ڰj��%�ޭ�L�X�d�/J?W׳�m]�[�U�=n<̀�){E���1�l�~���XN��-�|w\���J,B�ȝQT��mϿ)�4Z81d�5Ӆ����%�xZ~�Ӵ�&S;�:mF�i��H�ډ�qF5��I�n*VY+��L�s��ل1>��� 0��kw����1l�O�(#VTW �j5&��!�� ��Lub�5�H���37jd�qs3�oca��0��HU`��܏��/?�*�<O�zg���^H�N�g�e����漸�LX�_9�/a�%ޔQ6��HF];k��L���W�+l~�QI\�y�%Nrg��M�k�����4�6�8���v��ZZGI���-6;��u[��Q��s��p.0^fN��cJEw�p��gD��H�4mB�����±
�C�����eh�(���X$4�����c"��3�^�������R��\E4�����?r��nm�K���c;�v;y���M[6��{��I�%\!��M��rZ�����? .#yk�g�`c��T�W
n^Ժ�g��M���2����l������iBym�V.�)/	�V!�@La�0���n��b�}����a�z��:��6�D�O�(�������䍴�wb$����������0��1�V�U-�Xq�ݸ}�#VV��$����G��鸟��v�����!�?'ۼ�%�dj�7}�vM 	;\����|�נ�:b�h���[�|�:r�8 �j�C)�.\��>%���l�������뵯�� |�I���^��iB,�}�^n���+V3�q�������m��3.v��Ƣ�0�SVJ��yhѯQ�/��GM��
 ��T���˶s��p������({ƿp��wi�l� aFIV�~?�d�<K���u�*�XP�,��:�0`�[�]\8M���Q;��(�as� ����@��CΠݺ֛��y���'��k��U٭�E��ӆT�4K�p���zZ'vX�$�s�;K�tR	�,���:�C8��%�UNe9Tk�ڻ�.�5��=�:B}F
�Uiz����ʲ��̏�"Ϸ����x��a�s|Y��/6݄��ǅs2����N�7��]��`](�`A��Ŵo_]Vc��8�T��; ��+�1�O._5��F��]�ڡ�`ӓ��,���9�I���ӕM?uP ��y�3��6����hFvQ�0�^��\;�Ʊ�L��"�)ID� ��յޥ�Ui�j�vL.�q�ԯ���ԩ��ςz\#OR�їO�w��b𶐩 V�yD?28!	��S\����qd|�����Τ��ޑ�ٍ�;hܙ�����J�����8��>L������xE�Q�L�5�B?�H�>K�
]�E6���t@���؛�]�FV�]��3X�x��T0e$'�&�ui���.m�jʫ�)���F��	�!�@\A2�1$��1�큁8T�!@�8^����A�o�&���~�2���G�h� 18�r�}|ʪG�����^�H�h���Cr�Dj����l��Y8ښi���QP8( Qcu%�臄�0׷TM(� *WӜ&���C�G����]OlP��+���ȓ��[�����#ъ��Z��?ڞ����b'1�^�g�l�47��萾~8ΰ�{X����.���I��8n�r5�~f7r�o�i�r�R���.:R�1,E�[V��yhT�� �!W�'�u�`AOA���E��%&1(���l����O�O��'����x���$�2Zl�:ˮ�[�3�?~�y�*��|��JH��4���y�U��b�B�/��$��w�Ģ�6��Ɖ+���8��n&��헏^�^I��aEZ~M��,��n�}�y���b�֡U��y�o�4��i�����I)�Ex%��;��������ĝNu�l&P2ɍފ�a�	Z9����R4u���s� 4�� ��0UDPmXf�8�;����Ăg����s��hjIT�6	��A /���>S� щ�j�G�����]J'v*�Ѡ��Yx'Txo�[�lu�G��\�T���e�F{���#_����!� ���<'�KĽt[�4����1�)~)23f��֘,�2�3v���O/���m-�X>N��
g�s��ʡ#��"�<A��v�3-�1H��t x����Ot�kaT|s��L�׮�[j�����_�쏨%�;��'H��B¹�1p�# ���)�Ro��B�`.w�qb2�W��H��$�+p*`,�	%̵�kjo���G�q��{O�S�8_3�\i՚��"���lk��Ax�#������	����-�އi����N��ꪹ�3�2p;�i�����y���iO	�a�Z�O?M�t-;����b�$M����f��q��a�7-z�4������� �SEq�3-Ñ�6N��p(��4[�Eom�*~�3Չ�Wy�g��w�S e�MСy�e�?��������6�F0�Nʑ-�4��]������ V!-7w�u�J:�4��x\��8��ō�|��:xn^
�%�{F��"����(�cW+B']+����O (}����&-�:b9�'/��1[X)�r���f_�y8��+ �-���)�y���I�����5�9����b�"����4ZH=�!�k�Vb �`���P�"�쩕���-F�g�%�,�^"P7�b������E<B�\����Cl�K�5��g��N�W�B�C�)��Xhjȕ=;�q���0A��`~�����Vx��B�������YBr7O�@R=G�x*�/���2&���,6>�����=�F�L�����i+�H�9_>��u:�a|<pHVշ!�Y��`������GH�%�\�*tƨ[OO[X�}���G�H�?�,���<�%Ҷ��V5�in?b��+uD5�5L6�G�U�K�n�6y�FD����];������jӰr}��hJw	ş4N��Bf��L�M��b"�	ԩ���~��?�� E�Ȼ�@)�@�^���dM������1�D��Z����J��3��W�\�o0q�C�*�{'#!p
��&�s� _J�>E鸉p� �c#ʗ.>��Q9����W'�0x0����Foő��|�����w��&��n.�_0�+�������̴>4��U �*wkV��W�+�!,�QAY���
'z_꒳��`F����I/@̝j���@5ٍ͍��TeT�6h��>ӄ��;^��w��ͼ�z��Z� v���e�L�^'i�0��=(G-�熢y���E�dkE]���˝`�D2�z�z%\+��ph��g�%����i/=� �2��A�N9Cu��g��V��E�1�Ѥ���J)� �kk��q.��~�>�*�Z����E�0�"�1D���CHl�D�|�@w_��;r۱��J<WN���1�P]=�A������s�=.�d0��۱=j�-&T�q� _� ��T����<y��a�g�E4~����'��V�#ء��)S<�z�n ����f�2��1<O�'D����~9��HD�З�vO�v}U�T/OKU�Q��t�_���뗊�^��i��Sz�Q�xw������.�D��g��
���盨���Xfb�G_/��DKo��^B��Vwe�Z&k_]��ܴnp�S	{WX�JD�oV!��ލ�අY���[~9���6x��`l�,�a|~R���lH���4�h�q�4��s%b���޵]=R��\�6(�]S�� [�I8&���fCq-��Ł�����]�p5#2��V�KF���/ڙ�I��?�N�P��ߔ圣�%���h*���Q߳�U��(_ D~L6�:����*SHֳ�,�(�k*kK�l�?���r,r�#枪���.�\*<�T�����G��v'3tUC:^���d��u��2t�r�l�+�bz/r�X�jیm6)�x����c� �!�����v��T��>��ݱ�?l�a�~�~>���s��\6�ی�Q���#y�ßCՃ�a���f/�?���G�P3����i�3��C~�3Ɩ���r*�X��	����8�>1����O�_��!.��O���Pr��R� �;���稱/"��z���U)�"Δ�.���<t�I>�t��O�39�5����Bh'�%������}/�NCG5�8ԟ�U&��"T1e����ǁnXK��5���j/�"*�1��B"D�+K��ǁ�������@����n+d+>QjAG�H|�$P��5��2������ k_���SER�KA�J�?���4�~a��OQ@�FF��x�O+��N�����w)�VH�G*��57�EAJ;�a�g�?G-�d,� u�J�`�}���>~Y�R\�ŏ�tv��b�����;�{���!��'��Ϧܨd���~h.&�u^�����/cL �.���]�30��~���v���T_m�~72%�N�o�iz�����i�g1SI	`q����r�WL#�i�ZG"_`I�JQ�������M;�`���Ϩ$�oZ]8���岼�۵�5e�Q.ׇO�q���p�@�Eɜ}#c'�1 !�)��O�*P`���=�i�䐉_�/��sq	}ry��"����g�	QjSMށ56+�d���j�ؓB��׳+��.)M�����Ld�&��``��|cW��$�ՀQ`�(R�3�RTA�s�Y�E�u��JS$B���͉�É�ǩ���t#b%݊��LfrX� �G��M�L�]����F��&�s����p�m	�$��\�����|�`��l�vs�>)'XiD��]r }Ѱ��R���/R����b����L;ۤ��^=��~j��1�+�0`u4�I����G�� ��g%[�o��@��3�~���p3X%r	��;�q��,K�}��Ȑ ����o� ����P����Mǯh��r�!O�V����cK�V�l@l|0G5�:3Se�i���N�a,�	�]�m:D��g&�n,� �Y���<䛂�ϼ}F��o-�q�:P5�#f��R|ҷ���e����H|�>ܐ�az�^u	�b�n�	P�r��}q��+=�ƽ���1W���E�4=���(�dPX]�m�B����(�����kxܐ�*r����:YII�ۮ�������RV �}�Xنd�Լ�S~��ؔ���oK�}�'L�s��6�%]Q�������@��#�i��͇����8������Ny!��q��V׹����}e	�$-(� ��C�	cw��]��6�,{�/CMr؞�����G�ش�����e`���$[��̿w����-�y������������i�\xuK^�fŰř.c�r����a��Ӑ*���4�V0��۞O�J�pDT���1C�M`�u3���Ė��2(y��:��z�e}a�;%D�1`��a�˸��|���(>���z���!��"��eZ��C��d��zU�~�b�3nQ�i�l#�*��7���S�ٮ:դ��N�su�p��X��6ڑ��W��qKY><�"&�����	/NSHwJ��E���d�)� p)c�q�����AoÁ��Pt���('�q�,9xp�٪�ޒE������zt��4��u��x�0��.~ɴ4�1��^u�Q�z�vr�o'D���	��N؀֦7��Lmi���(���ʧwH����P�� N�?��/�����N{��%W��r����IKz�~!��?e�V��������x`;0.T����/�J�Y(Dv�kFV��n��x�˔[ܬ	�����Vd�=���l��L�Q����^�ad�k���D�x�}�2*B �Jv����SNO�3
�ؾ?�̹�ˇ��O��9�X���Xܐ���C59[���8I8^������� c;%�y�hC����u���MM9�� �J�K+���&B�·�$8rֳ*�#�u�l��,8�D3HZQ�\>Ysx��;6�ޚG�d�*������{�4sf�	��ɖn`?Q�`xH.��[�{3�t;.5B2�@�a�}b~�/BHkY~�^��&�X���7�3���&5������+������|�%à.ЙHx�c�����*o�_ٙ/���&	����1�(�`�.��,��1�������<E�~��w��C�G�OBł�u΍l�VW���n�OQ=�����VK_���;>O8i279�A) )�G$e�,�t3Tޥ�'�����g�42w?�_LQ�k��=Ƚ.f=�i������8�(���ݲY��3ҕ���D���j�kb��H�?�7Q�%-l��a>S���"锬�`9��C4?zΖp�U��gj�2���J�j�鹤�2���y�	�m���,��������ҕ��ftX��Z�~m������,鞳^�g[�W�Je��(5�ܹ�"��xv��gؒ9vANL:n}��!�#N t��u���3���|���M.k����^��S�U�?����-�,1F�e_�(�h�Fu�!��kF:ԓў���7`��b��4O����6�!�<�;����3�COTi���uy���i�׺y�=�Z_Y;��Oh��(��i�tA$����ԱJʌ�2�t�������a��-�E�D7���A�>�~��b��y��s����P���TB�ą�������ȫ�Y�"V{f�ްx�C��4����O���j[��Y�4J�iꌹB]�6g��Wc��@1\M�X�$�k�.�z~�������:IC-2'���Lv螑��D�T�����i�K�t�K�Zl��(v����Ci�*�&l����5T�����ͬt�_�r��4�A�Z�@���ys��[�s���UMtp�4��ju�7;���5�Y��Fo���~����<>�4
/�v���M�� �˾Y��t��:"x$�����F�\W����P`����<X��2�(����)��� er�Q��r�T�$ZЖF�S/*�� ��j���h"�����7���b�5������+ٛ
-�V��q��7��WCPBO\}�"k������$/��}� ϛ7�`�χ�7�A[��ݬ$$�����~�.C�WD]]|��a�^�ٗ��:���t���Iu �B���=�A��:[Yj������Ǚu�s��Y�Z�����/�T�C��I��QȲy+��ߣ� �Eq��蝉�*}���_�]?-g6���%\�Z�y���  Ӣ��%x�[�.�SK��;0c�� �ONΡ�
��j��#�
J%�*z���}��j�l�����$Z�vQVw9R�j��꺉
�'��/�B��!:�m����y+Q�9R�J�Nα�r���\`��(��K��ؑ�7g�od^&'�%����G�}�x�FM��ͬ>D֫�C�j��	c�}�lq�#\[������$ݗ����NM�����O�t� ��<��>1�[�3��Rsi��]���g>6ק����*�U�G��4c��k�n�k���D�JSiϼ��mϏ�H���f�FHQ)淨�*�.�t�F������?Jq�!=�Z�-���(O�L K�
�Oَ�,�W�<<L�`#��q'�f,t�S� ��0���b���B&`n��ɞ�����s�gI���R�1�}W&����ܴEj{H��y�B-�q�	ՠ��D�����J�[k~q��4�{恳�.�$�;+edJE5���女IZM�RIU8�w��y�Cvy}*(��؉ءC(>���p.m�#ѯ�N��jG���3�Fi��e䭿7M���#���!�o�C]m�UѾ���n�U��.g�M���F�1�:�uI�W��}��2�T㹁���޴�Y�����&�Ǘp�Hp���bh+���z�fvҳa��<�-r�2�u
�T*Kk�M<�Wxq59�QiT�(�R��
1�Ԟ�A�L#W�}6�_��R����������8����3��x� ��&qU��k{T�/�>%�%�I~���<�*���,2���Y�u�'�;�A<���C�rk���X�$m�
���moLj�.~L���w[�a�
��鍺��y�_#>'k��Æ�����"��kI�k�'�����`�����|�PP�5�������c,�y��
(��Ja��VV�R1���0�M��@��1��5<�;-�����pݪZc��q��X�h���$���Ʋ�����տ+V�KBQ�T(B�,*
�zz+�T��$�cc#��F��7c���Wd+�y愵��;�A\��"9��b�du>/�f��~?~�r>Sa�d{cĄ���q� !��S\�29YI�����]5܇�~@��x�W����~53:y؁d7yL+�)&��+�G%�˗v`�����'�y�j�R�����G�xF��fkQI�t`�{��X��Ό�y�3���z��C�>��s'cz�����Ո�+�a�k[��{xn�J�$1�q฻��(�^�� /*j�NL{�n�š��C��L�o�<j������X�
������op�!�8�O��hw���׷А{$\�i���āa�L8��;s.N3َXē덪��]��ĦE�Z�zꅚm�޿����=�y^��d�?gtUBFv��O���XcY+1OF1fi_��%�ސ!̾����(��a.<�}d����y�Hz��'��}&oT����V�;X.iN��B�A<��T�}ԑ��読�;�L�ɭj��ڴ�O�`��R�俥V%]��� ߡK���T�n$�0�1����ȋE��Ti��/@oڕXDZ�^�d���p�0���綢I�E�g(��33I#�����i�ǟC�����VXj�G�����*�0Q�b2�e�Ki�T0 ���"|��x�Y4g�?3;~�b`��V��\�Yd���ǩ�
�(H��_ÿq���t�M���<;h�P�;�L�?��$E��įB&T_�ƭ7�������O�`s�ܵ>B����Y�&t_��ԣ9u:5�a#p�<Zd�2֝"[�L�UH��.6>�h(�����kD��K<���?��)i����B�gҽ�q�������/�D�{�ǫ�7�Po��Boa�����ÿ;zNa�����_~�o
��􍅢���Pcr5�Wu3�z�OA��F��D�7��_�sG�rln� �� 3J䉱��e�	:���D���̇w����@\��%Q��Cn��p�E:�8�I:6#��Z�����&����U���c��@<n`rC�'��Jg�͜$�
!8gst��_�׿|��GE>YMk4�K�����T��چŜ��I�����0*�����������Ch�!S�� C�����MvÚ���3���N���3�[����*��\�C���}����6Oy^����H^hˠ��*�E_�$�����q;��t��k\`���o$7b	kF�<�4�G���a .�`�A+[��Lv�i;��.�������A�!��!āF�#)dv�1*�}�?�<`/���J͔"5J�*��U�R^���Ɍ�W�+zA�)�)����,���;	4�~A�kf'����p�����j�8n�^�i�p�<P�=���E���*�W(�sւH:�K���:��U6j���Mn1dݎ��&'�~����Xh�h6d/�-$e�|ͼ��	&k"��|��v��O�Y��qU���i~�`CR[���+��`�	/����[�+��Y�d.�����%�7,@睕��A���\���Ҹ���1b%�Iw5h��ȋ���ǃ�M��鴝ݯ�b���(�^RJ]F�}qW����+!��T��)~��'�&<�_t��6�����`H5J�An�����NN2��/�TǊ�>��M��n�����t��^:���T�1/�jp�'H�z�i9 �`�˯�p�eaΣ�%��}+�y$�&h�Ļ�� Z$n��M����͋��_�nn�e+����S
_[Fn���|'[��τ�ɔ0�V���Tӻ}Öf�AFm�Y326�VD�?�f����!��v$�h�ru�a�D�i��e��:I�x�G��\�B=	�O�T*ļ}sq_b.*}* ����BNRaӷ�]�K�˙w&��>��L�qQ�#/�@�+����^����|����,�54����KJ��/~_�F]i1R�Z�_���>c��E��1���p��wi����Y���)�AY,��ܠ��B�︷/L��j$`���&��������A[�of7h��{3�=�ht�'D����r���W�_x�_�ԭ��Yb�E�^����YIGw�����!���Q��!�_!�k!`���P����j��:"���\��U�@�n�>#ٜ���Y	���ysT���6��>9��h������%�'��i�	���=?��(;��5)a�,H="�H�	>\��7O@�Y���<#Ox�H\��m��|v�@1YQ���-	+������]7M2g������4I���RE�e��Y��as%3�S�}�8���Ck��eS�IC�T�.y5��O��͈��S{f�q�jI��o[��¢��ӥ�I��G5�Q�sq���:���d���xD������0���#[C�%'�B����+�����,�([$(�]�e2R�����;
�D��@���P��UUԝ���[6cѱ�O_5�Y�ul�wR�6�]2���f;�w�?���۵��Y����y�K���F��tn��R�8��|�l�W�3���S���yCn��A��nކF93��]1!(5�v���[	��9Ö\��1�,�gi����??.�i)����9�0Q�l��^1i���Y'�Ywǐ�u�D�Ɲ"t�H�K��F�MzM��R��o`�ʩ���G�,�1�]�S��+��Z���sKj�6��3��B7���Wj��2�p%��+�b]�ޜZu&��~7Z�Դ�ͳC}�����66BX�d�=�v�3���ݰN�|3��s��!�����$��
��~w�����P�'E�c �}PAPfʌ%�w��b�׽O�5� Ҏ��q��,�i��y��`��tX�/���A�2g����,�����D��zL��=_��������4;TѸM�l��&V������a཭K�)V��~ݰ:J� �
f���73��UM���m��v0*��iZ�hT?��ӊ\�}�y��h�!�('||b,��'�?�a/��mHy�z�O�����*��^t��nn�N���R�w�V"j�yPO�d��d-��b��b���!X!S,�P'|�1�t���~	6X��X=�y�/d'������\'���6~:��	�ǡ��*-�)�]7�p_��|I��7f�>
u-��9��[j�X,�J��$�;[�Xv�Gsu+(<�U
$% ��^�����@�y����׿(?���	�������`g)jb�LI�� V�y����!����'���a�֊�F���}/�J��ꢦg�� NN2��9���9pzT�0�"���n��ޘ��]L��t%=���o\3��"�LBݖM����%�qL�J� +p�f�I�dM�s�ȑ{yb#%���l��w]9|*]��8���?	l�Ux(�LN@�1*r	�;룻��2H
��e+�	�Syo�����ae��v�h�$�y��&��W�3!�z�ݻ��b߈yR^��Gb��t��݌�i�Q1Q�D��x��Pf��tG������֊`��&p��[Ιhu�tٔ_�́�Ll�����K�� W�Iy���"���B�T}���X�%{��^��O\�{ ׮�',�DI��w���9�dF����|AJ>�
oe3:�S��$ɳ�M�<�<u�
�tz��˷����b��$�cB-�gLH���(&����[H���P��:�b��3��9��N�F���Z�I�����PpN����r!�w�i�8�&ǗQ���	̀~F�<�D��w���9&�����O�@�O�9qJ��!����#CS<! �D+����"�9a JߟD��B�㓦i�x��L�gL���Ƌ5F|sّw�쳴.��U|��؄MhN/�u�Ǡ�[��x���嶀 >'T#�~�k���P+Z>j]��^�)���W�_H�R7h�a�
�·���%�C��Z|�T���W0�p�ےN�_w��/�-AM���s����{������k�m��q�bҶ�W�"����*^7��f����_�Z�y[�޲��Z�&�CĈ6�)�=H��~@��O/I���AiAD�Q�,��.#`K�l��]m��(��Mwd��A�a"^�i�9�{U27��b��A��Nfb�x�A:?]8��|yL��Lq�u����a�sGu����ܯK;M�����>x��:��'�H������N���`y��RC�I���{sǔ�D[a�b�E�*�H�VC3
)P�,Mɽ��ؑ� ���ΜuB�ܰ����Ay�[��vs����5Wq(A�)���cd,�I�oc_?��9
.u�c"2<M�Zl����.�k�jߛ�������M	wu5�ԋ!q4�'���-�^���,Q'���Ary��6ɫ��� (��3��I ��)�ts*"��ٺ�x�FKK�wu|���f�C������;�㜼�U1z2t?��jץ���yK�v��
bj�>գ�ԋbMM;$�G��B@l�AmOhG�Znxu�A�0j�ʗ4��Ţ��դ��d|�� �q��J`�&���fe[Ÿ}e���m�PlZM��f�����{Y�1N7o�2b�������ZtR�G~�b�<z�$;8e�=�ܬ6��H㺏C ��r��/v���>�#�V$/2�0�,���"ף/���6v��ze�
SC��W��ikm4�پ|���-pi����6��tl[���1RJ��c�|�^\ޱ0d1UN"yL�(�nK#��� ����Q���Z:�x�v���R������L�P���1�S���B��#G��Kg,���������|�ջ�+Vڑ�h�&�[eL9���8\-��lO��c���&�]�GR���ks�ǒMS'�|�u(� rzO;��]�X+�q:(@��D�C0�m��,aU����O�丮��,������͒M
�-�&"|U���P�U��HP��nc�k�/%���s�?R�p..�lS;����<4�ۣm�x��B�Q�kȄ��m=w�?E�2ZD���Q�cQ�����Y�~fUF8��`�Ek$���5�p�P���h�����`���	@��@������T��Z�C�mͯwa�k��y�2h�,u��c�- �4%�F�ʴgw�� Fh�A6��B�9��v���W晆�_���{�.RH��gs�W��EV'�f��ca�*! i�Q��#9�'�[��i���H%K�4h��=*������=��5��Hb`+0��<����7eV ����4F8�w�/h�$A ������E�X�p�M�&O��iHt䌸��`b�I�KK �B�pT��wz�db g<�8�II��y�k:f�E��!9�I0��'���Z�b����^e-3�)s몿mcY}�2�,���F~�h�G�4?���§���_�ʹ)���(�Jhm�!�5��D���A�Q-Uz�
��*B�\M��j-&� �RF��p[�W/��
��ݾ�N��L��)��|e:�1_�0��M��]_/��&��,ɤ�8���ڴw�=J����y-L�!��;��Qe�`��ֶ��ϵ�=H�0��De����,=YY���U.ٱ�R��OI"U57Y����cO����bse�
Q.�~��j�DkT�y��]{�\ж�o���#LZn_�%$9�b�D���q����Ƙ��ׇ�,��]-!��)`�^��ct'�f�"�f�E�^a`��b����u[�K9IK������w���R�&��D
."��AI�DR7��Ȃ��2��m������OI�𾒳,��w�g������t��e�j�o����&����Z1 BU���pφ���^m�A�
�]zfꦗ?r'���a�~i�mr�&_|V�\1�kl �[�N�~={DŁ�Z�;�e�-.&��ʰ��������k}CR�� 1Gl���6xЙ��3 @��(�;�f��<�6�N�[pg��Z���|�L����������M�"�?G��P�o�S6YV1��,Y�m0XR�R�:�o��Q��cpq�0&�0L�գ̘N���b��ǈ>*��84,1�����@_��vo�xA��#r�?y3�A�'s�r!�j��]�6��6�̇���;o��ℨ(�Fr�#e�.I�P�%�dע��P�}�\��TLɒ]j�����جț�#�@O*[&��&+��M;�������X�/'�����uz�T}�DK:u�>��]�p=��Pຮr6��+Gջ�d`��K'�Q�$JѰ���)����Yl��f�����~�b}�=�!T�y
|3_��#c���y��k0Z��Mw��J~|:��s������.��t�|+�*��a�1�Yi�*<W L`$�˘��zv�+���_C�;���_�V�����g����5L��ܔ����J�G8:��ҵ�-����Q�V�e@_���LQ���Y��og�r��ϦԢfM^;{l�(�9��S��ճ2�<�~V݈ѣ�A-��`Q��W���S%��=����GF�}�ҥ����pE��3-��u^E�7X%,X1����X�wu,�.�v�j��e�-z�H5���<DZ�,Y�y����"\����A�a~�~�oԶ�.g��pڅH�WX�����C���s�.%��Ou�1z�U����4u�w�����V��A��C4��B"�e��^�]��u֤�[%.UC��_e��H摂I,�绸� I[n�f@a����>�i��ϔ���qT3K-Q.K��k��mMJT7�u�ʟ�5�F�*�H��,��H{�C�9����~�C�fe<���܍iX��$O��\�Ȓ����g��v˲�٨A��P�n{�bD?<q��w�xJjAoa��r60��J��Z��#.�Cj̩\&T�_i��b�H�B:8������97D��I�d,���g���yݣԗt�����X_iト)��r��q�S'gFdP53����n�M��Hi%<ƐL.�hh�5qe�3�{+�񛫎Y��T4I$���#��M�7 I�[3=��E<�5����?�l `H��&
ϯJs�c2��9lV�8�'�~�s���a��6�6���e�Oq����Q�N��_@�[���/W�(� ���6��|+Y՜N`G��KB��r
��R�+'2#WpDG_���_	�)���b��͂���T#�d�/A6ь"޶|	�(kn�@��7�7,�:�~t�A�H������-���0jI����%�ԝkf��y�f�P3Q����r&*�b.�8�l鹧)�7�eZQ����/��y���7�l�}�l\N�16L,J6?����4��tv0�Aa(\Z~���w��l2�_�m�82�^`y0�j��&_S��f����\��.�".wn68|��;%��r��4��"I�LV?nl�f�U���T]Ə)�0M'�K;OĠ´�hel���#ܹ���T�U������z���|	�I=���"����4˱ehqaQ�un��k�J)�,>4�g�b��Y�	�]�chF�{���CP��H�N����i�7�������c4 4��`Gqu�)�\��O� 1�~@̮���4i��HK
���zkS������<U�T���s�:��i[������:�P�?��j7`vo\�
ߧ*2��J���N��0�j[��l%P8j��XA�m����rd��_��HԈ�kr�v�&Bu5��'���)S��Gd�� �6Z�� r�K:HD�E؊%��2�G��� Z_�?��~1�u��/O`g���TWۉ�u���_f{Z(hR�+>������Qֿ�ăBk�֯#e�ry�����]�$C;=��B��E,Ԝ(VT���WBs��W�uVG��Xg����/=9��a}�D�4��,�f.����{�8�P�k(}��x�g���|�M5��A��#�k��'����D�HS�O��^s��&t#�;�1�Ewʪq�`�S�)�RU���dK0F>�+��^D�(Z����O+KXIЫ�� �J��Q�E7�;����6^F<���At�:k�)��)J;:a�k�,rv�cw�y;ǿuIip���n���|��F��d����f�ux/�ձ<C]�T�T�	q�@��G�^���:g	 �:���=�e�v����1��c�8D���C���湂P��59CԲ�>�c�L�A�/ǜ�U-T��1� k�w���:ZJ�l����=d�d3���T��:��S���vl�UC���U�&���=��m��Ȩ
�rJ{C�9�I��7�2���g��1��i_	��m1 ���~>x��~��"�R2�B��p_�߆�c�l�)�����I�9��WіH�mL�d^��2�W	��Q�D��fR	���<ˍ�ʡ��oz2��8<EJ�H��p�&�kO�g��C�*+�
!��Zm�����M�`�Ӷ�86�Ly]WZY���1aXWU�L���B�� =�d ��]L���Qbp�͝�1`0㴳��\���h�k��*M4��2:��zc�����I�*:D}�)�~6�j<�-\�on�?�=��`�O��>'4�}ۮ@�R��ʧu	��4O�y���Ǌn�q"��/�X-4<3-,j�GO��1�1|�[�:��aWA������or�nvVР�(��A����mMa-D�A�j|Ƥ8���4T�Y�2���b-}�*	*� `@h�E��[��'�r�8%+��y:D;������B=���P'�D�W��kT�T��-���m �~w1$(�μ��ksOֿ��L�é_$N<�_���?}dE�ݟ�_�4 @���Y�ھx�ݣ����N�׼g�����8�(n�ԩ�a��-�@��Ya���~�%�M��`�w�<�$��Z$�рH���n?q7'��oB�G���v����av�߲�=��r>DyyJFD[��`��."�3�$�0���2�H`���ț�N7p��oI�V೪k�9D�2>v !4j���(�
JK���sc'cT�#�Rb�����	�X�)u3�Is��Wkd�rd��V`B�����p�PiY X0��(*���A:�i�ג�	�|:>�̻ � �R��s�};3K���$l�������M �w}�5Ě���n]�+����
��� �X
L��"h��/��p�E�+W�߄m�,X�9I+7�8}�|��thڵ�4��FI����X1i�y�����<L؀d� ���6�-#�ĺ}��>����ʘg��0I��G�e7��<��ZR���#�IOc����&|byp��g8 ٸ~sc7�d�w����bd�5���LH�L�c�`����>�*��KF�^����XT����H�F������<k���)�tq�8�\�Er4?��r��$~�Ԃ�tbKqb�T1,Y���F��e
���뒰�7��.$�feg���y�������
"RW�i����%A\���G��e�х6D�Ip�mC��b{�o�g�bzT��3���;�e���*��%k�"na8�s��6��,��p�ZVHR��G%E_�����D2���%���x0��)o,Wn6�W;��~����VL=�&D�à��쭢��ߓ�;38���+�.5�����ծ$��<*[G��֧HfX�Q~:ېX��|P�~��K8�w3�X�I�p�����v���;�e� *�n����G2MO�`��^�|R�ҽ0�2���XU4���#5p��z�-�������L�j��t�fy��X�W.B�o&@�?�)�le#c4H�_�U��)�%|���W0�[�k/W��D%�~��#A^#1�>V4*��;&��c��m�{�u*Wfd����#��:�ۍJ��'7[���)��D�Q	Ey�:Q%(֍�P�W����k��~v�xSӮ�>N��A�*ب.A��xs!2�F.���2���c�w?�ր2��s~���E�%j=��n��E�6��%_��X!����<�J��t�-�E��a[��D����~΍n$(�7�E�����W;t�3�:��$aT�w��� ��iB�*1G��CK�/�/�B�/��Z�_���4���0�G�D�#�倘e�	�z���t�K8y
��=d�{D*�b����(��C��L5�&J����8�H�Ѩ�Q��C8m?�7���ɾ�`LX���W -?7��;�����[Ӵe�S�*��͚����Nہ;��Ȏ�gr��d��^,C���4Bd�y��K`<��t܁˖�2B}�u�nҬeo��H�꧑�z<��T���(bOo�a �>;(����+2�fɱ�&hY�T�2J��f���>��ߧ-��)�Aҥ3��$I��9DN���5F�IȞo��8�� L��N�ʏ-p�];=��������Gy�33��2��=&?~��;�L2�(�68�8S9l8�)w�@#�!ғ3�O�W�Z(�́ȧ��)�0#�J��e��S��:;�R+�=F�E�Q��mc�9`�dC0ji_���2��Aڵ��\�.W���Z�~���������e�Z��/m��Nz"�	 ޫ�vlj2K���D�ߢUQ;���B�e;Q�\�����T��'.�W7���"1~^��e��Q	W3w�����ş���+�(~-S�VJ������s��э9o")m��e�xpCK'�7$�C�+=���P��9�M��z�"�IZv�����'�_�Fb=�*d]�d��ORޞ,G�)��W�������c�Ζ����Tz� '��s��a΄/,�]�5�V2E�\���k�a�`��·4�K������O�1O
���t-�"�2U	-�e����6�0��8���R�~� �\�w@b/X��Q�U�%$�D���^���=R���Vc]��Yimx,6b���I�ج{�T��v܌L����I�� �g�Dփ����,�KV�ݬ�X�U�$�o&S��|�b�� 4,��ӏU�h��ڌXp!x
wS*�!
��<�[�L�Eȝ����G0�&Ea
;����2Fo��}����xVZ4��h�����F��Յww���o�ʣ�<�Dȕ���A㛏��	-���9D6Kk�ܻb��!S�ÉǞvo6Q����)��s�g���!ю��
{���|701��k½\;�A݉���{���[ϰ��|�X�c�ps)G"NX^� Y�-����'z���^e��`����!�}u)\�c��C�`�C�����{8�z���,�6��8�ޒ��@�_�{���T�� �����,��6����� �����S��9`���,+/q�k��G�T��dO�$������̻s����D����*@�ɝ� m��T� ��]ά��@Lj���Rƈ������������Uf�^y��E TgU�@��Iᵂ#�]��G�pDh��������Ta������K�Q��|�~Q���da��(��`�^-�(LWA�"'ze��?����~���G�N���1�$��>�|󝿉9-���l��F*Џ��7�F;�b�6#vY��R�� ��T6�H
E�����
���3��m�`Ց�6�ق
��P�F��С^�\�R�A&	�l�0�TIm������C�q�	�Z�1�ڹJ6Sd�
���N���~��D��sߨ����fR8��	ZԻ�����8�&5�ůq
|)U��v4 �rj�܂�j-�x8���QI�� ��i�GƁo�w[�F�����SO�/�����ma��{U�	�u�x��f}�P�^"�bXJ�Fd5/w)bk=��d"^��/��_n`��f�}ȁjN����J���io�W��£UPRn.�qjMV0}������ �!�V���TS��_; �,�N��r�h�4ؑ�pBScnKA;�tUZNXU����0� e��#Y*���Y_1��l��_�e��7�u �Jj �CSZ�x%V\�z�>�X��HէF^5�
G���	3�Xok� ��"&Έ�~Z�K���}2~�Q&h�7 у7"���f�c?w?�݉R�
` ��I�Ӳ|� G����ST/�� ��]T�C����1��'!;��od=�f�����4���
����y85�k�)��l�8p�)a��c7�͟�)�lT��E<��z�	y�[^�;��k(��}.�4I���}�����B�5�O�k�+��כ�%d@	��%ʶ��� �4�P��r� *aZ��K,,%��l3Z��<�I
l��x���N[���+��=C�=�n�?�� r��.Z�3�i�Y��H;H<������ۓ�m��������[DK�,P���ك�Po{�O��TAo�_K��I������� �/�6v<� [���jC�0���.��h�^턌i�6"_�P�z3�廨fgNA��{Û�����%��|J<`"�7G��x�EF,nb#w����s�5l�d�S_�)��P��(�zj2��C�:�Q�*��e*����E���I��<���� ۆ=݈q�45��8*�j�<v��R�(9P@s���ʡ���]4jZDxy]��u����w3a�Д�W�֕
�#����·��@�\>��e�C����,dK�¢b����1]:ү�vz��X��*]("*�v{=�v����&���ƋY-/@��L�gI�w}�%��娳���-�z����܏�`����D�w�6_����Gt��K����
@Wꭞ~_�,�u-��s��A�C��SH]\�����d���f��Ig����|����Y�`g�a��^�`Ű��!uhlg(2@
lӛ���5��	Jyn*�C��A��iz�K8�9O�W�eǤK+��4}��a�_���r����[�/��!<V���/��}��c�Ƞ�̕�sϯ��FiE�z���`"k�a����h����T����l~�)!y��R��s�?˽�|<��]�8e�两r�Wn3`�ʤiw�
a@� ���(�3�&��@4�����qX:�f��b��S	��A���d'�8E�*�>(�]NaCj�=R�-[�����I�)�����ܪ�r�q]lVh[��Vm��jt����a/Z�t��w38�85�Wy6܅�����{��|=#'�����
R��=n�n@fZ��.y7��m�۪��ԩ!������]�g��]k�~���5������ vp��H&`����g�*�:��\�&TT�ޟ��=ťf�B���Q>��6-�q�\�X�d���jaj�Jaꃠߟ����L�i�+��(�|�h����V	A�C�[킱\kb�j�'w�lj��rwcb������*���RO�r8�j�=.i'���=/ЂC��H�оu�Y���4iΑ��^�2n��)��P�m�gM�Ydǡ�S�4ބ-����݂3$Ҋ:6G�'�&�zW��Tt���HC�Ѫ�jWr~�a���?��Gǝ�'L؃ѝ*���D3~�ݷO�ت6��3SRԂU�BQ�����~�iWm0�	����i:ow�S��W��3�Eǘ?�[6c~���:��h�1���~���gmXxȔ���h��;��uP�z?�����N��J��,�X�4su�t��j2�q�)�FؓP��ٻ}�la�j�-[�=�E�)�x�?�A����RJ�x����|���w?(�T��CBc���N�x��$��L��;t����z4�� $��ײ���Y��	��2��!�:��sm��]S֑8��W(�+���i���!�,"�����;A(�0(��*��Ȯ�9�<����&�3S�S���"�?K�?>Uz���d'��,���S���n����z����#p�v�Q�S:0'�MU[)%=L%�c{���~�$�&�EEE˝��Q���)�G�E���{�i^$~u�j�N6������h�����}���K $Xw���D�Q#������� ���R{!���%/�;�Qw"�C3S��{���N��f@L�7J�ȁ��6����Ҝ�UԦ_n5e8e�AC�l�v���`���]~���ÊP�{Rx�
�/_e��p�wj���5��<j���F��x�0%��1gA�<����!���[Sjt��8>����2�����FӎbO�$
�m����9��G$E^1p%���x���I;��;<4Rh�� ��4�(�EN�l ��B����kpNb�b�Ey<�YE�p�x�b�[�n>�����o��I�_�zrn���D��5���!O�Iz�a�|6�hxj���b-�̽��X�)S�;��T�W�P�����Z@�Ӟ���['巣򷇿�=�9�T�d�3��&�3z�:ӣ7%nm�%�Y:����)C����*oXwM
L�3��a�E�vv�=�IyT�tCp#�k��������L���u�0���~�}T��I`Z:\�x�q�l����#�nن7����čxGO��C�/��d��\�%�A��$,�[3�r�~O���8QU��M����#�9�3ܿ
l�f���K.��V1��SIB���K��ag�E�%���l]�u>f�x���z���&������4���<:�N0��>7'��F�.�%L�iB'8&l�-�h� �(��޼"���Fޯ�!��S���qh��(�g�?#�$�Zcmd\.��a��/#�RQ�^G Op^���������J�F�MH�Ӽ�#O��cAձ&0i	
@���$<6�ýG4�#Jɂ
����A3�r%_$8�PVz�7��%ԩ�Į@�9���N�n��#��$D����99�:n/���Z-��_XN���T��b��_�prt���d�f��P�#J�,���֮��T� �ڮ��9͍�T���}6Ss/Z7��aLO��d,�cAaV8�]2�B/�̐]�pVi/{��W{�h��� 4�	1��]��#����a�f�e"[��fc��`�"��g�X���9���#~�䷰���E�6,a�����^�֎3��s!����K����hp�K$BWP�b(�Z ?u��;�D7���cV�-�Eqx���d�������%��;�#����q�����b�+L�:�d���4K���.^�x�S2�Ofa����`��4R���Ͽ�ˁѾs���D�{�V�q<����)��I	qF��Fl�N�M��t9�A��QP�sd��@	`�J�y�6�/bn>��a�0rM^��aS���'���z�v6�\I6����zeŶ8�G�5�Ė.����Ȍ�Gm	��ּb��ޛr��/�Lٿ��&���{t$�����4�>~#$���* '�Nf����#��c3&[狯Ř�/���t�%_�2EgS��q���S�'��\(�k�P?N<������_�
�������yIo���,b���\�ÑD���fX���/����R�A�P��+wV�R�5F��ű7/�t퇁2?�߲�ǳ��W���TC�/[�!�ꋸBS��>Y**B"�(-����ۄ��EMsC#��wU�Te�",���'*=�0e����{���^��ze�o��Y<-���\��!��h,��"�l���$%qgR��ɧ�i��L4���ߺ�ԕ7>���z������~�|v�%�B"}2n�K��ؓ�)YX� ?EB.�j2铿.���ɐm޲��V��)�G��%b��!��nJ�=5v|��Qy��E�6����$�v?K�Re�g<[_絋�c�F�%���	���g d��r�F����|�g�?�"��@�n<\H�K�G�H�Ј��U�f�����1k{>3��%RI9)�,�].>�;[�h^H��=�����V��j�;�x!6^��c�����*O>5����f�_CX��$�R�e����^6�����6�Zm&{�3'��f��_�d���w��:��qEH�l ����yf��~/���Pe���34�D;�9���.���\�'=0PB#��0E�Q�y"J��`�>��M��_s/G)��� j}�oO,��P~��?��8da�o�����ټ+ _ld�I������m�)�D�e��h ����#./ r�.�cׁiK:_�NY���^����@�
�B�u�DD	�+�� ��#%�D�����#�h�5����xS9����_+���< Y�����i���p�!�9�bKW�J4���3$��s([�˴:`Z2���~"M������wQT��\�C*;�zw�s��(}��QB��Afq��ĉ�j�i����stVg�+/�쩍QK��3�B��;)z�Rb�')��MsR5��e!+7m&2�_>�	$�b!J�glY[-.Q��徎C��-.��\;�`��٩�(�}$���åƽ�tӊq�����+᫹��#�5j�n�c��-%��V��u��+�v�n��z�0�!�z������`E���&y}�}�v�/�Ed-�J@�D�Pk2�y��֩�����]�n�"�I3�\6�G@}.�J���fG���O:�N0�I 
�~>��C���|E)pN��mZ�~��8N�T�T�\�?�3xLլD/���������N]ݤ��GT�5��Sp�sN8�5��8$�k��h��΀t
��m���`̙ƍ��ӂJr��6'�>LԘ��̊��GR���ԙE���G�8k4!*r�9E���Au\*A��&��y�HK���<�5|��AS���m�$6�x��<KJfj#�B�8�K�]F��(+��U����&H��ɭ;�(�T:p:�e$�Z�Q,�l6�>GT���Ұ����>pm�1_��8�)��2����b�NJ�c�\7�zƾvU/"L�uM�-:mGS�([�Z�׬�fϚ�/�~�����#�b��T�O�_�Q��Ph�"Q%�2����957��}��k@*$��zq����_���h	�~�B���)��v�Ɋ4�:e��2]�������,:;�f��Đ���~�lt��k�(ҟ��#�Q���:
1Xڟ�a��gJɹ�b��}Po��Ig�L?�v�%��n���2��[�H��8̿�oS��q	�� ��j�i�u���̋�G3���%s�Z�}�����5��7�t���;�o�!X����KD} ��f�3MN�D���A�l�PΠb�a��/��^�=%���A���q8�aa�?��b�f\�I��}��l�x�9����>&�>*���Wɣo"L����H���>Y����ŀ*�	�?.��=���˟ITo�Bjo�}��Y
MJ} mB+2B�g�G���8�@�}yRF����\qg�t����
�m6������Z��4w�j�o�W�j���C�0�)��]I{�?�L�>p�:���A�t�X�r�\�����"��u�)p�Oh��2;����v�5f��xk�,�{HJ�{�x��$(��f���r߲v�Qx{��t�lJm����,���,��'OT6r֩�]��Vr�2��K��c�${�r�s�M�\�����_W�sW|�5��8hרd��ȹշ�X�i�L�����Ky�yɻ�f���F�!RN��8˸u�)fie0�!'���=t�J��/Ҵ�ceX�/N��Ϝ��:eD��qǻ�v>�i�Xq �o��};ʷ7�R�|lt���k�:w��Vi*L��x,�D܆�L��չ�e ���@��^��o�־𨯴,����B���]������B�p��,%y�1��o'��f��K��S�*��_H2U��K�� 9C��|�U6,u��4�l�h�U��*�v���� j�j:A'��n���z�P�h�:��v������՝�\	G�FV�L�p�L9?ӫ�5�&(n��j=�Ǐ@��ܑ�'���@0]+?����X���u.�O�I�=i�	i�X��@�VTj~hv��4A�Ӓ�$��_������ݽ�㚇;�������-��)�z/�B�X��c�����$Ts��~t�\��̾�!-@t���R��vna��C{\�K������+�
��	��Lǥ��������&Z��-�I>���B�<�'K����������P{��b�{�G���ZbN�m��	3kI���U��/�x^�sP�(��s=��C"��t����T%/��+& ��.r &�y����1�m���џ�HH�H�����j�\��Q�Ȯ=釁��Ap�>D����vc����1�Q%����0�e�.�:?�lc �<F}oH��t���v�t0��W%^2�,�3�ί`f��9i�@������愦N������Va����n��k��5�l�|l4����f��f������:2�u�t�$`��_!��/iI*���Hq�I`۲ߊ �F�b�C45I�d����5$ybm_
��L������w?�[)g��6���O=�����m��E�������}��dX�KzH�L��:DE+M
��*�-�w��@��;���!��BH�fWuv�wե�*k��i.�~N���/	��Bs�[������qip�/��UMl��aD��$mQ�p\]�Y�K~Z�c�= ��4��W� G��O0�M��T���h#)�ڈ�p��}'M9��O�r%h tC�5�����$o[5P�hm�'�y��V�R���Bb���A�$��gE�ˋ���%��f���#�S��'��$�'�j3Fe��,�����=���gx��1���qc�\�u�XA4�m���
&�v�N_ž�Ү	U���/v���얅ޜ���C�Gv,~r�a�V$ 8b�D]��Y�$&)Im�Q��S��+C��[�9l�	kR5�r���`�a��lǢ�q�YOHݺu
��� �U��J9n��e���'�I��~�ŉ(y�Nb����ԧ��K�� �/'�!��b��aR�_����u��P��b��vh��ud��\F=����@���⡽͹�����G+3L�:u~A�s��׼>���b,�\�M�J����H�6j9�������0\����	&J8%@E�cB%Gt�e�O���b5[����Z�a�����
2'~�:TsO�nP�"�X�jNy;����9I�Yc{��K�姺�8���*
/;���+I�<��4�-�u;�nJ�=�;�v}��]�\�N�n\�M�rP�ju=f20�qቲ<`.�ǈ2���Kz����fʓlRL�͊�ZrsT@��������H�̆���_;�f^�����IUL��TrY�P},*�+��R�F��z��,���ޒ�\6R�}G�&6����H�n��H'%���Q��0/��G��D}̓��/��>���j*��<ʧ$�ɵ����AT�\f�����P��2��:N�|�4��m�����'6��u��G���u��Z���C����%"�T��X{�C{��J���e{�M� ��V���&�#~Γx�qt�H�_n����E���LM~�V1�6�J�;;;p��ˎ	���i�<���'�k����e�+H0�I���p-�P�U�����~�ō,#W��
!��	�MQ��>}g���>����W�F��c�� ����Q
�����@6��w;9������O�2Z��V�1��� �?���� �����#���l҅�g����S���!}@���l�~���ʈ��3�1��9���?-�m�ui���I/檡�O	�LnAp�ޝ �Nt��KS�Z@��������[/NTi�z�����>���L�  jy�דW^g��eM(��s�PQ�@��Lz]��]$ȏ��������χ�|9l�O���}�bvSv�է����J�ܥ�6��_�`�
p��ɯE�w��M�z�$V����E�0�h���ܚ�3�]�J^�'�%Z�b"y�ė�|A��!J�B|�5h�7�q�H>G�ˢo*��a��x/w�WZ�N�ge!�|�v���5�&���uu�����A�o���7[�?��������M�XG��{��^,q$��秕�.(ָ�柉��>|�ZΎ0�_����d/�t�"��u����Y�[�����ժ��!�J�{0�T����H���E(�1?�嚯���j�S�$E\N��`B�F,�s��i�8己��-��o�\���B��q�U���J��{���cu��5g��������M��������4;�z��GK��}�80hZ�*Z�z+�z5���D�%�e�R�:��.�?��C�����S��%��9/2Ҝ��v�It�B$ ݘ��"(E�s�&� ��m�2���o4&��j!H�Y4/+�؄�T\�/���8��^�6�1�Vi\�z{.���}[b}���&��[��f���m��?(�2��XV��?P,��ӾDN���cSaVD;�Jo	@tB/k8��;�;uܜ��a󘫌�ѡ��4��R� ���];�����=�.�M}��I)˧i#r����H��3���C����C�U�����C���af�"r��
��gN!���N��u,?�b�T�ʗWm�R�E;OP.�=%\�;@�:k��}�-��Z������;������B�'�$����ڴ�/Ⱦ"����{�e���-~W�����ݰ�3O�-<d(<�u(���t�'���Js�g��.��љ��56k���ׯL�!1�s�"���$J�`6�P���se� Ff�V���U�#ƅ�������8��.)��n���+حn^���fWg������Ƭ	��Θ�v,k{�o�z���4��u'�'hAPz�hɼ���v�%~1��A�#i��K9ං���L ��[�a�T��x5ڤ?�;x�s�C#Y@����Uy��Y�c�Z��U��k.��i��C��щo�0��HW���l�{��[���k��P�(����<��L�Y��0ƉN�����c��q?�lR�D�Zܲ/l-���\A�jbLIE�5a�s�7��8*���M9�p�49�9�I�'�i�e$r��)�/�k_����T��I�؍��o6p>���I8��B���&aQ���F�Ev9욍g[=?g��)s����{�p�`Q3rt��Nڊ:Q�QJ�c�)���R��@cϞ�2x ~*j��&VUK��ze�N^�aOu�G��Kd�t��Z�<f�����A�5$���ba�מ:���o�Sw_v�$P_���t�cm�B.gV@5[���L�iF�ÎS̀W��qX>�˙Oe��>x�G^q0m@�a`(���Q��
�m�z�I�%�X��>j�d)�M֛c��P>F�i0ބYQf���M���U��:G:H�y����������,R� k	��I�قl��9����P9���x���r,R\j��)�1��gH1+�����h�T��o��j��5�~tJ����3U�5�l���Y�6��|Ȉ����x��!K:y��G�B9�j��ݾ�>jҘ4��H�u�5*� �Tj��cXg���=��K��R*Q�@K�n3���l;f��胄ֽ�Oo�5�{�bO��˼2(*s��b��9��nN�o#^j��f֝�?x�ᩌ��d��|2'���ғg�S�G���^���=���«pw��?	Ӥ\�������?A�����WD��L�^ʬ�[�bJ	�b����Y��j�Ci&U����R�?,9~��P�i�S��Y��<U�D� o��	�!R�pe��t�L�43i����ƺ�9��C��ZL�`c��a�_QR/"�NLz����ݾz�hQ�A�75-5:�3}|��jaMg�%IA�7�΅q���y�d[p~T�I['������⊐?8�6z�Q��E��G�r����h���e��i���|id��g��N�D��W���i�g�e�d֎?;J�
"
�B�L9��ﵭ�N�d8y�D��i�3���F�q��������bvW���c1+�=�6�9��k3�jZg�ӧ��LÑ��2�Is�����	���_��Y��K���_��7����F���6�Ģ��//۫�~�p�R�&�й�����?�𴜯b;����>����J�Ac8gU�76uLcO�Z5�/��~u�`LܷNmG��Ds�48&^$�:�{{s�v[hn�[տ����Vk��iS/ ���ҽ��1.|�(����3#���ϗV����ųc�A�Z�"�,;�j� �64����vg����['�Y!�[�I��N
�{���lj����?E���|_�4���+�_��¬��,g�#*�Ʌ,��0�%�G��q�3�ӱ*��8��7���Cu�RY��)�(�6�_�ׯ�j���"�0�*D'/%��V3�����A��;��)� �z���MeZ��TXx�6����X��l�|F�;'r�C��c#�'N^�J�C��M�~��5A磆[0͵�H��l�4�����@��Hg�EL�k�LX�gA�𷅗MԖ�ʋQ�7�Խ�Mmo�x�!�?�X��j���<C�;0��)������l	1�m���*�y9Ҳ+�Z���>w��~�m�y��L��AM�pi1�#)�����C�;�2���89�s7��B�{@���=&$	l����ѝ��/\y�{�n�L�P��nuH~�}��K*E�Il[��%�]rd�?�6Q�g
��?Yg��B������)7���1S6dYư{:q���<ڑ���<ɉ�An��!E���H�p�ª�M�勅
s,$@6^���R��ۑd�U��U�E��J]�gӞ�v������(�e�������}`�ӐC��<��B5��������l?�5kl��q��?�^Q�V���G���0���c����B"��Z|7a�nJ�f�KW1n,4dJ��w�gy\�V� ��]yҁ�u?�%�c��&[��R0�E���X���|q�.FbG�3�b�4XV!��������'��m�ut��_뒒�b���Ć7�:py����2��O�	�(�
bI��Y����3�B�p<�;��_Zv����=�Unܟ��#Y��B��b�/Ðg8˦�	��U��;.U: ����t���9'�TDҏ�Jga�Vj��a��@q;�����bJ�}�KL�پgY�X�.�8��<�(��,؈4��:Z�`٧t+F�2n���|%I���Ԝhr����~`�#/)'��5�{3�z�c��Ta�D{��>��n	��(��j-y@���w��]կT�W5��aLeJ�$JA�["Jbڨ�AK�᧿��R��_�.g�G���η��f9}�R��O���a�ie􀯠��Q�դ�l܍��r)4>3�y� ��rZ���9Suo �[j�������mR�f|m?���>�7�=;WQc�?��Jp%@�FWuS�.y���
T/y7#��I4��0N�E��&D[�
o�m�>z�>	'�g��H>�̋^�j<�9xH��"T$9X�c)�_��(x�R��H�U��H�Ůޱ�>����v������o�����b���
l�"�ݔlV'�ύt�A��$\>Z�Ur$�n0��O��� ژ��^�������?h��C��E&a�h�U���u4�\�Lɷ
<�T��Q�R�DZԖ&��S�7@��S��n`<�'m���Y�}�������3&9p�0ʡѕ�V�#6�D�3q6�B�y��Y@�S1| f�xs0{Œ�l��$�b�@rtI��p�&�y�ܼ�EZ$�h,k#��9)2�SH��J��N�
WP�wF�R�߯���9'���4��Q���Jc9�$a��z|c�����L8�__���a��On(��|��t0��*l�J�{��8i��bM��5���&�G��s�,���Ra��_3����aO�VB�����;��5!ɰ�!�yS��z��XS��eނ���m	�*���m:�0>������;ҳE'%P�S�o=SN1��x�1��d5�/yӺn��jo��m����/6��XiI��+: u���B�i�:mN�4��|�S��bϪ���1̫ů�J�
J�Mn6.�8XeY
i�Q���lF��A�	��yQ)Y��[�'�9cd���W�>h��dk£M�Ďn�c)���~���t��i�oyDb�qA�
���<���w�Pڽ�P�/�;R���~��?�o�E�d����e��@�>]���1�-X�k~9�Y����c6n=:�
��Sp~�8�]��2L�!9<�q �2R��d#�w��y����Z��}ڴ�	�w�2)jӞs���l��������$�%#hNp����үK�:��|��^�!�v3�+t���2�����6��x�'��M�Mӗ�s�����Hf�Wo1��2�b?�?�<��G�S `�2�1�/]L�F��J���T�o�Y,�+=�b��s���y5�Iͤb��À
��q��x�Ao-��Ul=5$%�IIj)@���]R|�/����<�=j��y�s�t��|q�8�����|���	�~NgX�Q_�+��iݮ�Y���b*���57��*"�1|�~����TJ:�z��O��I��������{�}�����q�`�ѵH���}`f��h��5��,�-�n����8���*��Ka��l��s���Jk�,��u���ղ��<�EMhP�e��_l	��"�e0z����U��hV2��u��U�����G'dyrH�����׎�2�O���f��j~��+�w!�R ��2b�eCnM����*�W�o'�#�����j��v�����a�J\(۵����^Ʒ@Z,t�;��Ȳ����o�,��#����Q���h�p��� Ò��y�JPs3�U�;�ϖ��k�R(��Pz��G ���:А�?�������(����Cs��cO��m*����drYp����ފu&�l�-�����D?�`������r��ܥ��S5����1��[��k̢�k�J��	q����R1���sF������q3{��K�L���U��x �$:~Z
��'B�r�:g)0��d׆aq�u;N�pӘ�r'�~�3��]fJ[�#T��+UyR�+*�<��a�c,wc�wx�#Rb.�3C�,֩jh�����t� ���hN[�zQ׋�**��)w�����5b����^�1�^��pL}�����,�GQ��X���
i��j�|O�2�gֳ��|ĮisA�6���iؠO�LJ����߭*�ldP%m�j+�9��/��:#[*���J
ګY�c25ަ$׹�I��Pй���ᶳko3w��Msޗ�Q�fE����۠�Hd�"�w�<�X	�+�'�e���L��~�L�q���h=��4[*�`������¬��O�:�R�@���Y}`��x����c�R�$~�jMJ��x,��˜C��B�*�έ4DG�t���w4��b;߂�Ϙs������F�4��C[���cB�z=��_��t*��%�
c�SZkά��{օ%k�8�v+L��8R��zB�ir��`��G�(�/</3j�ik"Z4K�ޖz�z�	^��:��������N�9]|�0���:����x=1��T�_34X��]mjO �\�9�����A�ٛ�UY�f���� �F[X��=�,uN:���qE��2�̲���,���*׾GK�K1��Tcq���R���&�綸�f�}d^�1�?�)�l���;��^��;�3Ɵ2�� ��2���WiΐJ�Ӣ�	�aV6vU�t��<Y�]�)�;]j*��V���r�`�"2��s�ľ��Gb�[��Ư��{nw��h�`8���F�^D���~zbQN��k��@L�8�/@���Eo�xP[L�ů��w}?4�7�0x���q�0A$�"x]58.��6m��C^�$C�I��Xc��
8��b4zV�q�D����C���Ȏ:
=<�؈~<�毅�>���,=g.1� �i��I�M�4��Ǵ��}�V�,�A����/A�#"0��+r��nE
��s*���� 9�ԥz�F�JM���U'�GvП��G6l�/���nD��,������2��Y��/}�O�q�\,)���Q� 5��dL��G%q��D�U�AL՟�3�|�r���\��>�6z��W��C1�(9	��lS?Q���$=���\�}iwߜ�$
���-�F��!/ݎϝ]�kr�j���v>�4:�OJ���w�
������:<)k�: ��c���f|�����eW���m��<�%�W�ʢO��L�OI��ȝy��D<��s>S�RT1gK������^4�v���wi$j�Is���]�l�}i�-�r(._�=�5�a�A��`- ��K� �u�NC��` ߫rM��	DB�/���kI�=��D�5�M�r�,��{_NsO�ۖ�b
��[��d2Wt�H���ѾX��OD�FO\S5k�v�M���NXGU�|<��d]���Y^�CI]v���Q�bvO�+V�|��3�,j��r��*��`�1W�ύ���}��W-d f���Y��n��@�N�NF���x4����ե�Ӎy�QC�����ƽZah!;���F�\5��#{WH��ꂭn��äG�sUϿ���
 ?'��	�M|���Ԙ�J�A�!��VS�D��L�$��ş)#i���M͞��P�W ��3�"$�< �yȨy�8_�թL��ԃ��/��ݪ��ă��c�v���nz�����^�d.�z�+%RC�����X�e���;~_�e~p��s5[93́	xĔ1~����S!"pm��7�E!c@V_7�7�<�I��7�wEM�9��s�کxM7�����6���W
�.j�bu�	���➨�3��S��������p�X#�6��T����ޱ��p�/�T��b�s?8�6��Ĭ	20���T��	�O �O�h#<^�gHq�|�mڒ43�lW�]Na�E���M뛉֔�=�L�ec��?*a,āe�  �E2�I&�/2b�w����M&��m���*QC7���L�%|ڶTGNVT�22���B����W���#�ײtU�y'&&�����C&��:;_�λ��&��iEE��j�B2����)e��&9�&���f����)�3���Em�,��T���0�L���T�҅��6.��X9[n����=�#W�d�����Q�0+��q�Bc�~|�w9w����Uz/�� W���)PmEj�|7���0�b7�� ���$7�^|g�N}���b�"s�ɛ�ӭ s�A���8��I1�r3�a���a/���6��E�e�yFJ�z�^�MK1\DK|fu%����+D`)�Z���zRw��&@���y��'�h	!!R�8˱ ��o��3��¹���y$!�����P�Fɉ�y�R�v��R(Zl���1�E,~	D�ܺe%���oN�.E�Q�'''{��(�䌀u�	_f�}C	Q�WJ��[�/!$3�ꩡrm7Y�Z��˯�c�Z��\8	�V��%��V,�"T����et$���e�RK��*�Z��y�����)��� n��R��V?�@P�_r���?���Ա�yqju��8�@�aHl" z��ra�>j>�3���8 ��	 (��Nh��Γds,����	�%'>9�u�}��iS��wr�������%�ft1�}�l�^T,�~A,��BΕ���b�ZN�?� S���/k���x�qw�+?�3){Vo(�7Y?ى���������4w�I�u2Ӷn��r���v�D��� �c���;RSb����yU_�ysT�N��ӱ+��bY:��2����֤P)>(�t��)#$�K�6w���q�eM<��!ǂos��*A]�D(����a�_��ܤ(L�2�#̎i;v��J�ˉs�ӯ.��>�)��Ekj:��۽4�|��qDM�ʄ�"�R�d�tc]p_����*b5qP#��o�Y�>��!\r���{�"ݳ�_��ز}��G�i���dt1���2��.B�^�0o��x��+��1`�ݔ��jgv��cNw����5b���c%�ICݣ@,N�DUy�ҵ�@'�B�T����}�Ԫz���{���]&�Mx���@W]�3�g���su�j�۫��.��M����1�[()s���]�7�0�eR���"账q�J�����߅�؎��'��������1�"�y���KԪ����c�`weƍF*έqL�>�n7��<-�tJ5���u-jD�.Z}@���}�>�2em��)�1��RRqA����j'�L󾔌C���"p]J"�/�A��jl^aT�NQ�}KJ��9s �\\"�%<�O>~f��V�l�jƢ�����cĎ	+���i�סF�=�W�׌ǡ %�C�Nѷp)e��l���]@L��C��l����yМ��4!KL�Ԃh���Z�Ić��%X7V�� &)3�54+���҅OB�����đa#���r�Q�	��چt��+�Q�'hP�����/2_88h��U���a��;����T;?/pp��M4�h�,d���捶+��0P1�V'0b����+-�p�����+"�7eJy�/C9_��U%�.͊G���,I*�k+�6y�Z4֤����PZ.�G���dG���vC���<w��%<l�&�4������"�gp��%�T@��Aw���Ӻ��v0l�|��0ӄ}/�H���D�� [�%����S�դh�TC3>�NT,3��i�T���4
�i��[������RijȐ';�9|�	�@��-�\�u�eu�d��j3@HK�>sIՇ՟6��HXX[�S$���&�6�Aҩ�p,p7�|�B|fn�~��E������I<����L�r��Z���JX)W�3%E�(�P�������_u���-��8[�(k��d<����%�+�q�M�p�L~4ҚpwL���
�@�X�O�f��A�),_Չ��#�$�{ʪ�q������#�K-�2���3m���Ψ@�ǎVY�}972�|���(`��r.6\J�t-�Z]���Y'r�q�B����,w�~ ���}&�D�}X�$�&�V�l�z��)O0��ό���w��u螡���E�p����E�o�8w�w�&�{R�:��<ȗ���x�M*�W����j�A/�p�3���E+F����0MYP|
�Ǥ����p*"�#��]N��t�r- Wpi�˃p�!�B~"�:-�M)z"�\�3+��bT�X��[�9Z�f��D��}B�37�^�D�#�`�u�td�K�������$VT�e�b�Ҳ���~N>w�z��)޽�)R�­\e���a��c��Z�"�"^?�I#C���|��n�tq���$z���1GՋpqȘq�j���Q_Z�z�?�Ϛc�!lK�;�g�w��Zi�}�}�G����N.�`��ct���{Z��_Ah���"��y<�D�7��o���P��;�
\SjUK� eh+���W�z@����]���)r�U���S���SO9�3]����k���4En6���+(P��W=��8����r6�����a5�t�ZW��T �yv��3"9A�;���ae�qz�iB�ycX}���mt�Œw��b+iΎ�2)���
7�:m_�5�D:�M��矤�WX�
u�ɐrea�}8	8��;a�}?D �㖷��ŋ����s2�n<��"V���nio��#���ԏ�g�6���0I��a�|�r��X��OªXp� t�k�^`X��=O��G��V�2L�l��0�<^�*�i��ҡ� !D�?���i�㕗��"���(����*�[o]�����r�#�`	t�c����a��\�_#���&���&%n �5�fT��l^�c�����
`3Z��Nh`�IH=3C�����Q���$�O���Fa�U�,�tI�0hYf���@�Gv�D�{�%�'z�����7�f�I�}�H����j����oӠ|,����z_Z6S���_~�[�j4��4�!�ֱ���K������,��啥Eі�ˌUCo}e*�x�f�\|��&cB��qՂOը@ܭ�RLF�BL��\?�������#�IV��Բ�lPh���sj�ܘ�.*i׽:\���H}�<�	�O>M<�%,�{K��~D���	�Z�c>�,����_F'��]�K���=z|�<���h3l6�ɸ�t���b�MR�� �;��g+f�xb�ۗ|4ȣŜ�+����M�!���i�����)�Zm��ksLY8+u���	�F�JSs$��K�p��j�·��Äx��"��t�K���|���|0:9<��2n�-����Ǹˠ(��I�m��Ñh,ʑ������tU��ީS�o��<��(-'��$�����B��pY�t'���>�j��4��U-}�׫l��~H�M���阖�pf����F�MUa�bE�RL�VL���&2��k�Z-A�4��	���K{�%�U�r���]�!�����j�;�:`"�K��w/g�#H"eB��S��u����Z����Q��+�u̇�|���ű�WO��̇
���g�Ų�B��`����^���ǛC�(��x7ƣu:F���KZY4~�_#��]� @�sa�%Z{rxw�T���aYx�z�l��~pw��q��ث��[P���V��[��)�DG�H��fa�P����˅�Y�^	X��*¾�Vb�v3���~�p����{�Z1k�ͦ�[,$2$O&��p҃?M�f;>#�	���)}�����s�2V�vO�g��"�0���B��v��8���N�������S��8���+&�&�z����U�4��7 a��a����	�ť/���Y�D�&G%�[B��cd?Xnˬ�^�(��b{i���\������ *�2k����#d78km��.��S��a����@�T��h	���K�,S
��6��4��F�\��L{� k�$�����'z�@!�; ��w�U	ьB�/�
���%!mq �V���k�/V���i�̴�Ǫ.���Z��Ti��@��d&��9�l۷���g�t2���e�� ��� ��NRV sju�9�c��Sd�^u?b����%���;a��������)�l��N^��)�(��|RR�s�{�S�@��tS�y$�#���)��A��g�\���cW�j�z�[6h���V6�p5V�JB�u*�J�K%U��>c�tn��qǶ����}^�m޵7�Uq&��
�$ժl�9{�����������miB�	Y��<�Q=��1aT��c1kãt�����xd�T倝G)��?m>�(�����\��4�`s��Fb��(�`/�}��W�Ƣ�k�Y8U��M���)zꪂ߳^x����p�� �{�����B��|��q��z�k�18d���%��SV.��y�ck�*g�#(����־���<���v�&nk(`4��0G�q�Z�2���$K��N�h:�&�ǫb՛��̂��$�nkV9uV��;�jk��J�hP1�����B]��g1}4�t>��Ͳ�9xT�uq)�gX$�*�n"g,m�I�J{����Q�����=EI2+>#w���QJ���I*gh��X��B︢�o��+�6� `pKF�S�2��[bV!����TX�ci��aU�\y�2�j+��;����]�!j|Լ�� og����pA0�O��Jmrׅ9<
�¼�'���sZ�C,P�~�9��'��Vyα�̼7���_lZS�!qfbQJ%G�6��'Ұ[��$.�P�s[���?��;m�W�w��	�8y"����r��Y�<�OJ^�Ԣ�3����}x������8%�4T�(NS��u6���x�E��'��_�mH�܀�
��iQ��\Zhɇ����`�۰/�������p%�0E�����݄鏄�Fz��>�Տh����2�@���:U��+�B�j}i= 2s���XW�v8�_ȸ��yb�v%//f�D�t�`�L}s1�Ri���z0(�̷�����}�eՙ� ��YǴƬ	U�BNX����<%�s�[��9����;3�p}�A���&`B�ؑ�5��c�N�(���8u�A#�Dk9(����Ņ��`ZU��i�aQ���`S0|{{({��$��@H\�Bc5Ŝ�p��}�qQ�K�x���M�+˙�|�ӕc���F@U��8��h��o�7�l3�2�.J7�*�L��h@:�l�ʅ{�����,΀���!Bܦ 	4I
yн]� ,m��a�m�R���ĥ���[�v�I$L����=��O�$F��Q|c���_��� ]����![_k�E.�i0��J2d8r����y��Up�+ЖJ#����by�r��W�B�7\�I�؍�o��.L�CP�\�#N��D'��	�:q���N��{[N�h��f+3��c/$3x�a�P��	K��}�7�ǝ�^���,7�|��<<nO��<�2�%J ?��8^b�D@�k���D&j�����#_@>�j���� L)�S�l!ó�B�%�X˧t�F�Υ��-���r�Υ�)�[jI�v�h�";0�x��W�� @��Ưl���L?�M����N@(�������3�c�o���tI�n:�c��S)I�/�g[�˪&�մ����d��0��3�[LE	
�>�v�ȿ�l��HH�W��ZCp�v�i�x�3lzs��l#���xX�E���P79��� r;A��o�c���ɠ'�$;ǳ�r��rc�%E��bh(��LN�8a ����?6xiJ|uB-1H��?.gj�5�- ��l~n���m���JT�XXLp��Hiom�~[��~�>��e�J71Y����'?,ԗ̂�Y��G:g�zʔ(���e~2�5X��؉S6��l���W���n�?�|Iltλ
��SB*W�'[O�CY �hU
�ӌ�`D�����W��U��g[�y}� n�z �)x�T�'T���p#�S�Τ���c��+q~�N�|�'�)�o8�	�=&��l�0Q��:��`Oل�����^��է�~G�5k~��3ig��Wa�>�����,U5�<S<��t��t���Y���%��O�{�Ԍ�X�����&R�bR4#�aVJ�|2�OᔤV+�?:��5'�B�	�I̋�$�Ƣ�#?�)�<
jF&�_.s�����8'�8�w�ۯ!)�|�Z�E��jP/��6�|����s"��7�Wq������\�}�n� cA��h�Q#K�x�*��<wq����B��BO����ìcH��7#�}=Ar�{���>r�y�}��HQ���:!X��VlR3���]~���-]<D)z�^;�'5CYnd�#Ua��9n=.�xڧW~�R41*��-<@.�z:Rۇ�'�wt�#�o�1�ߝ|$�xM���p̵��2|E��QT�MMϾh�+��C<�s���p��s�gs�]����q=�J�\K�ŹH�J�۱�G��`0��Is��-Dk�1X;+�i�C\���E ��+>L��-)� .�f~TlV�6������l��=��?�&��^@��YZ#�?�����t��5-c���R��V���#��lC<�������l�sw ���gڶ����§_�^�iq/.��d�"��4����O��w�t�S� I�_��g"M��%�N֣0M�q��WCۢ3�����M�4gn��M�N>��=#��/ gd4��=�({7�~����i��G��WL NVu����72�����6�C��k������GE��jD��������Z�d����&�'�6��l:cق���c<}�,�j���/g�����boߧ͂09xΪ�`����S����JDq�}�M���;dZ�'����jj9����4��YR��!�Y#��
;[8�����+�{���Kd`���r-X�:��8��Ӏ=��Zu���"V��|��m�oĮ���_Ú���q'o��̹[��xW�T��3�"Q��� Yv����22V,%�u�ȋћ����q-��|�5f���ئ�wV�����D j�D�coܝ�"���)gsc`��:����U���%��a�B�
/���;���	Qώ/���J��X(/:�b�D�a�Tf�D�/�F[�@,vkm_0@��5GȈu�iw��kb�;G�c���@���� ��K~�AQt�<��@H�:��Y����=W�p-ެZ�T��З7��z��Dڴ׶�K6�#"�R�#vTIb5�jX���'�S�����#<�S��o��Ok�������v��i���F&/=݁��jrn74y\�`�{-�E�$?r ����N �̬�ʜx4A�P'u��N�^���v^p١����_j��hεW���L��R�GD�<��?K�53�(�< s�B�p`�`<r�L	�FU�G�*A�99��g3F�ܧ�|kO�!!����Pў�]2�f����F�+ F8]Q��1��N�����o��M�T_E�lD&Ǘ�FI��  ���s?n�<9�N�'��7{��z�2��ֶ�p�]�N&�[�s87����)#m�ABK�L	:pE�'~��m0�Xm�fk�o��̀o��Է��_�@�*�����@~��.����`'�틇9��z�m�x\5�g̐�b_]����w_
��F	��ԉ���?�3[~ݝD`/�~���_�66L�}���8Q�t�=@7��[�J,��@���KD𩧏��
�B�dZZEɝ��N Z�[S�೸pIx��|_���&�n���;ƀx`��]�Sf��V1r�r3�lv13i\�̆�/�����\�N����;cf��*���'��T!0b��G��~�"T�3Hg�B�.��4�8m}ʡ�6;
�����lZ�;H1�/uu�)��K{�Dy;�T�L���c�5�m���k�o�l>��#қ�W5�(a�����*(/�w�6EÅ���j�D�nt�뿿�YՐ�<W�F���C����IMb��y��J��R�2K1��ЧLr!A�:�ޡa}�8>"8���|�^�dbr��՛�c-u �O��7�c�7��t���k&��',z�b��|3@��Lby���3)WV���"��˵#	i)GXW��D����!G]�����*`�(�+�q� Y|��B��*p���٨�l>Fs -���.�*�!L_��f�����M���!IMB�-�6���l��I��#��A*��b�ce9Uڤ�Pjm��p��k/>���]�6h�HzHS�c�)�{)����ɫmc��e�~%�!�$n�����
{ShG�	{����
G� �&(���1��b��1''��\��>�����<=�$Ao�������ě�-,�2.z0����'�z#J��Y�D+��׊S۟�;�]�L���_��^�� REkQ~���Xr���-�I���z�W��!Y��k�;��E��Q���
��ȃK#��:У5�f7���X�l�\;2	Ð����F�;�~����v��zW�@�"Dʗ]Ύ� ��5����2��d��u�,��itd�����(�l��Ȱ��7EV�s�{�l6��?��'Tq�`&�DK�]C�3:w�,�����F�[GA�M�|����c�D�W�f��ۡҖδc,tۤ� 5K��R??�t�ݰף]gX|��K's���B�R<l�e�����7y�j��`����^z��`���N%�XI�	����,y�%���ԋ�$�`��\ҶJ{/�s*�G�M��0Xc,�'R���}2F�E�Mw�2"�6a42�L��?�c.D���)���e��j��g�Ј7id{�k�G��|W�&H�����K_�:�- 6+8܅s��A�T��j=F�ʶ��V����Hn��q���^1.}�aq�.�{���`�������v�O�]���7 �>�v錛���T�iD�E�(6�)]�����>	yRe��I M�̍@��K=��Y��ib�����_�Q>4Y��G#�Gq�4I˜'�����z������	�{3�@C��MpM1�����X�:����^SVU�V�Q?ҙj��
�!���������S����ֱ�P�U�.����0G��=�N�d_rxU��a�'pI4s�"�];.d���x�ٰ{�5h�B�ƕ�N��/a���X���Ii��b�h��\���i(@���)K��7�Z�*�ѿn��ǔ��w�ߜa�V"÷a���l���GGX$K�=���Km��B�#R�Ƞ����$ſN� �w��9h��5s=?�/B��&#�IM����l�!�f�V���/�'�doQ���ݘ'�ZN�V�s��$�6��Ç�#W7̌�91I���`۾����{�������1N	�aiU��N�u�*ϩ�d�Wգ��tR�����T�-����,g<W���w���FL�1�3pN�D����I:',Z0n�oi��7���.�~��W��ঘr��5NI�3���?X�<%_%��	�����s�f<��,��)Uc-	���Xܶ��t���:@ze��VE ����:��s@����p��rf��R�k�)�w)
/�"�<�ɟH���Tr.�D\�I;���;�'���E�Ǽ�{�z_k���K��pfL��Y��j�H#�Nk��`k�������>��cV{�0�O� v9F�</�F��υ% $�d��lH���|�]㰥o'
'�y;�6'?�}^�I욨 �`�n����  �L3�	_����z���-�Ϙ"'�|����q�����ǳ���Em�2&J�,a߂�I����C�e1�g2������m㓑�Y�AV�^�b_��Tj�6#h���(O��C����ƕ����I�K%n%޺m��4�~/7�5灷7��%r{D|�uǐx#�Uf�p��eʬ%�b=`�g����0R�S��2O��j��+Ȩ�?�Ni7�z��.����`	��j�@�O���*'��82��˩��zHF�Q1����L͇̄_n���K�
��Z�G�ڒj"�y�-���[vگ��L{�o��Mο��%���I���P���`(�6w��l�s}#��9�0uv��|@�����B�y��{��Xy[iT��r(S�t��w>�Oʯ���=�)�U�W���L1`O뾟C �E
�m��6 i���+�7���}�W��jmT��q�!E�-�O���[��lA��[}�o��RH��+��m�\�7�#�:�6Y�ǔ /�v�s��U������MA�#�k�Gr���s�JXӋߤ����z�4�p��<���\$�[Z����������X�{�-�#��ד�H�\k<>��Q��ʟ< �
l9ip��&n�h�	�)��������eGJ�.�O{�i*�����_a>*�qJ�68�+��.!��m�͈,���A�қU�	��ɽG��M$)��?a��é�VfȰ�ͨ/�d��ZK�>���E���m�A���̧��ݓP���F$�b#'�,�]�K�"�"	����S��
�2aey�������, �[_
�Q��Ez%�Ncc����gR�o�;��v�C@p���	�=_]��%�w��u��95�~H�����n3ٮ�3�x[6}z:G� C"�����9,�<'�P3����яJ�Bg`̦HW����l��]�Lb�2~^s�iŹ�&%Sn#2(gz�2����1��X[��n��i�g #��8ۣj�*]S&�n�G�7�gy3����Q�̵6i�\�9/x+8�0��t��.�r��hc푍�s4��e�7���e$H��#����2h��!D:��[������� a�YGl���Dٍj��_g��봱��uW`z�xi)r�������C���O��#�-
6�-�2��	��� �Y�LY�6!�+�Tn�ʭk���AfF(����r9�E�$�W���i��4�]�����6��j���Z�b����m���lyj�Z���/B�	�i�u>�*b3~0��/"v�3�mn﫽�:!^�q�x�	K� ��b��1��/2��#'yv������}�9���lϙ���ϻ�����o�;Bo�GF�]Y�,a�[� ��a��VLw^ܪ�-0��BR�#'O���;��4p8e=����:إ������Z���̊�A���c��Z���@WۋzMLi�m���'Uk5NSr*մ�}�3�2��������\Z������k+՟�e�O9�zG����c��!�D��)t���c�� �>w;�X��8�qd@���/�g!�x
r�~:��"���� �ң���q����
1��W�x@(�-d�ʦH��)�@G�^Ԑ�"u���V§JC���0=8NV���}���}|r��}*z|���0�����HE�0�0�wݛ�,���e� �
!�m���X���nΥ7zy�		`�Ѥ�YH��_��=�8���� Ӓ��� 5*����(��k#�1���L����mq�YfȖ�ZB� ��C�9�+$ĒJ�����wd�N���j��:�x�gPn�2V�f���%�p�>��^+|�Wo|~�p�h����h �V�Y��8�5��8�cnГ�ʰU̯m��q����hI��+�E�%`����Ƨ@��tĊ���������й?�zg\�ϛ[R�P��������'������[�F�	;�3�OH�ؠz��	Uc���q�z���<ӚƁ� 	l�Xsl,:&J���>��<��/�AI�3)u������%��"���QK3��+�ns�i5���;6��.�LkP��ƒ��(�>��C1zs�е���� K���l���H//_�]v�BZ_%E2~C&o��Q��"}���¢�&��S�UOz�3kj(5*�͵1�5�0r�.9#�&|G���6)�k�����:0z��&&G��{e���ͦd\1Q�5�DWm�9���A�և�G��Ъ���8)gZ>$
"*��3�=姄4np!=+��m�f�~�����-�ÎI�/�+X��-�z)�KAz���(~�C+�8
6We�oL0�SA��+MP��x`=�A������@�%R��{�H�v�9�D\	�m��M ���0Vȁr��Z�[��W�<I,UQJ�^�nk7w<����Ga�-�{X�9�񾤻HƒR?[4�)���Z@uIN�j��z�&�'b�G�o�%)!ޥ!|�BuO 1ƒ�L��D��#��RۤkM�\����?;����}o	������q�H�{�@h���iU�S8���U��-��jJt�Wf��n�({T�!�،�U5|� ��Wlks��u ݅� �DT�/���O�gG�Ѯ�}�ƭ�(e�}�ڭt�_x��?� Q	D2Ũ�1}]�Y`j�,��c�K�9Gfi����ג86��Z�Y�0�Z�wa�ls�;�o�@�[F�*��rL�}�{��(��1V~�`,.A�Z����ų�e����>��/��� �Qz�I����x�8$,h�1�ra��|x�D��1��|���x�3�2#4^A�)0�ϐa����V5V���M_�>���\\�k�Hԭ�鋈��}��ѭ�ܯ�2Ѷi���` K�	�b��G|�q�v3;R�Γ˯adpx����G��������m���SHV@����
�b8D��D!�F�f����	�n�[V1O!��%���v�6��HɄ���8�S\�U�b��Y���p=�ڷ���nj�:�׺���>�1Ɉ'T��ֺ᷌����ՍOE,[ÂY��	�~"�h��ec<���r���H�N �hBe�����S����X�������!��x�![��qͻ3I? �RSWG��Е�{GZf�Qo���;���=��&��Cl���PQmZQ<]%�	�㛚͡���1�_�?���Fq��`nLKI#l>� �̤
�1{��p_�7��,TO���RV��Ǣ�n�K���9�V��F�. �!`R���@5L��hA�oT� �f�K��Y�L�@7�,�S#ћ�J}M�y���V��d�_==�,�\qU�&�'��~�Kj�wE��k?m�L���Ul-=[����t���ڷ�zw�@p,��o��
5[nc�'`E�"g��}Y�Z&���Z�Zy[�kC�T��d��S8��@��Ud�`�4�;\8�Z5����=P:����ql��i�mٻ�׷R�h��:���G�\#AL%P*)��O���0?~fz��}��8������˖K�H|�'&H�~F���4�p�=�q��)LTL�ק���R���Q5�M�M8���e(��)��3��##}������&q�#���!ý���W�ΩU7�8��0T�޸{�O=���!l�����|LH�2�l򿩪Z�Xf�ggH�����Lj�����Y8�V������'nf��u2#��ׯ!�����ā�X�w�(x@e;`� �"';%PNV��B�I"�՜<+�(�G����Q�E�~ݐ7,�q̤�I�����Y$ �Y�n�"{��F-���|ȕ֖#dX�#ED��9���������2�5��_�Z��SO�q�d^
r�<���h�5a�p�z�^��]�9��@�TѠ4��.�9�ˊ��qH�	o^8Me[�*Ag�U�=�"�A�>0���1M*��~�����`���佁L@�Jc��/^gXq�H+�ݝ�)n�¾L�c>%�T���,z�]�� � T��6�j��~F|ÛkV��}����JZSrM�JZR������uS�	��_��5��O�w�ϫ*��l��t�	x�ū9\^K��h4z*��YI�	�P��PW
E䫀��!-�f��߁��;Z}f���G�i�ˮ�@r曵���g�fU�r�{g[��9{Ʈu�wo,\�9�_O��u�MԵNi�W���%��A��k^���.��vXCs�����#���,��E�R�� ��Õ1�	-a�ˎ���#��lGA�\�#A��3��t1ΧB�l�;�",�,��6��!�`L5�����>U1�llF�I�V�2q$�
&'����7�}��F�{�wI��5�����}>�&O� B����v!c�V��X���Q��]FL�#��˕�T��(:���Q��=�!���8?0@=iH��7���XP�t8#���/�D���L�}�T��������!Ul<qט�m9E1A��v4�d=�����4�6̛�9wp^"n	�=�&�ݟ>�������CX��J�/���S���	��Ķ��4Ph��4q�|~�s�Z���Ĝ"�e����e�[J���R`w��3 )��~����K��$�1��)� �<�jPg���zE�� Z�8�l�S�Ud~�ބr�y��ǧ(h�*,n���VG�b��V��Ż�2�۾����?���j;���l��Z��^i33�rht�8�ۖ)8S7��_�ĺ��[�̝8�GGf�f�}�:�W� &�V3%�S�"��k�4�fa��Q-E��*dGt1�=�3ҲS�,kj��ahdIPӲd�jE��c���^�1� �u&��m�&b�c |dݜ��������"/f������0W\���N`�;�3�͘VW�C�vH|s5F.�F>	'TԞ�	C$�}���D�J���#ݻ�5���y4�����k�d,lZ���4��xD��ղw�B!1R��W�1����3Y.���o�}�mm]��SM0r�BMκ��u�ұ8=g�1*�ΰ�ư����G� )��v�� �cu8)�3 �����N}-3��D����������u���銏�I\W�QH?�8r(~��^(�4t�'ɵ}����]ɧ��3B������iia�R�	eZ�6sS�O�*�go�]6D�0�32ZFӵ5ތ��,E;�[���q��.Ɏ/���<*��q��9�J������ה�`�Q���Ϟ��鏊��NI�!�\`��*���rB���
�Ù8�X_3�L�G8�ܦR�S(����hq�x"�q"�gʐ$��J[c���q%�n�s�HK�C�HUs�]�>�)f���CH��\]�c��oJ�n�
ea�}D�1�oR�C9�g�Z�^��s,f~8k7ƍ�����DȽɢ���?Ŕ�V���pr��},�Ҵ��>R3Qԋ�;fc#<�
�)R�g�ckw
�uЏ$O�Qp����'J���i���[8�^�T0�a#�ۨ�ڡw��4h�GD�j���9�5`�;o���_it���a���������δ��s(�[9?��Q/a:L%c��A&YRI��JK�Õ!H����v���.���rS�GB
��!�&���}XM$�X�7v�7>�&@��uSa�(N��y�e<� q�.)"g�آķ Ⲥi\�4+Y�N7>jйL�̐�QY�����z{�!s��PWd�#8d�{u �J(�GEM��u���`�T�T��;�*!�����:�PC��o*�K;�bax]��U�j�;�	�gJ���Vj9���?�P�%En�*�6c�_�k��\��Rr?��Em���Ph��[�a�=iS\4����/��N��+��s��A#���/8pi�u2m׼�,ݕ�|�,��P� B�$%eR1���ؠ��j`F ��{A,+M.ɚ�=wI���"�0�T{���1�
+p+����d&�O��?��\OV �#4�'_�L'a1@F���\�ǨES�G�k�5t�
��l�ݚ����ϩj�Qm5��/�������.b�EcJ�~��u��}]/�ϓܸ��>�"F�4׼	��&~�0�s`�:Q'h�3�`^�(�i|bBZ������9�Bq���#�M.7����^�S�v4~�t�q�����EI����{��ֶ�fy3y�~�Zl0}>��'��5��#+�(MI�,x$��7��@��j�{�[�u	=�`�S}6O@�m%k�.`Qe!�m2MU��N,j.�'�[�3j��2O��z}B��u���X������|LfHu�?H��7 ���~�r�oB�P��n�}Y'�σPwM|�l.��*��*D ��FذD$���4/�o��^τP�{�+�.�r`���-X��ҍG�K<	:� ��1��OKh._F�<c�
�k��H��&�zD���te��I1A�}5�Ԝ��"	Y�XQA�J�z�A��I�,�U4@�G���T����g�yL��	\�@ëH���3�0�6ġc�_}a6��x�p���+f'�g�Y[��P��Y�
6}z/˧j�"d#꜄�r�aRŔ@&F?c������f�k������t!��k½�I$L��%��#� 5�%pY�7I ��_�*�꫺��-p����Ǌ��,��0�>���i�
i��/PC;��u ���k�y��:��\�݂��;b��Z�n̑İ�'m��ڱ����J�O���� k;�$�ʖd,��q��B@�y
���k�"�P�V4�ơ
��	�Dlj+	P4Ƞ�rM%��h1r�N�i���2��iR體�5�R�{u
�04fR����W�Q�#�bv�S[��x)T���s@)γLB�l�?df@�xҜ���S`��Oī�m��;X��/"�/�;ٯs?&��Q�|*��Qn�����%!�=�Z��o��U4��)'�J�.jipQ6��x�5*�(����+� f��z� ��1��F�(���
���a��JX%�?�1&������]���։-��glD"!6c��l�|� f�����[���ܨ�J7�0���&]�$eŷ#!�����L�R���~L���������ih�m�md*ҷi��{�v����/�",���#��:k�KŞ��Z�=�_���L��M��R�_WĦ���[u���!�Dg�h�mZ���K�߈CJ]�j�;�T���k��͸_q���T��=�|K�%��z�mnr�K+�B�'|4���6|[�*����ۈ����4I0�0��˛0�kﳖ8E�����G��)<떭�+��"��������W�`�I��'qB����$�[�ٴ��:�/ 5l�@Ch-I�ۋ���e���C���%��d�z3�\�*C#���9N2lnf���Klh����p/�~��p�r|��y��I@g!�_Ƭb�S�1�(I~,q��"� �ȿ`8o�_yK���1��c��N�q^X���)�H��On堁0�$�bS��`��z���c��^������J#v-�T��H��CJ�z,�������Ѱ��K2�V����M��-mO�����Rg��7]�0H���{�$C_Q���R2:�2����!J�|��a��y�((��ѳA�S��f�[?��[�Rz98��?�Ï4�F�3����'PJ1)�)p�4�wuT��!rC6RkحSr��h^W�1T�����|��=��q�9n��DC�;]Z�.�����s��:�H��q{g�@�oC�C�~��l�Jg`uK���WF��N�a�!��b��ɏx�d�J�W��I�l���V�tr��@���Ey����+u2uւBIy�%����Ԁ^<s(��bl�����ށ�a޲B��.�1K��]�O�/��&Qпz��Ѩ��|�7�l�� `z�x�hҀ}Cc:3P�Ђ�rpy�Υ��wBW���TI��h�M	�횬9ѺH<�#%nQ���up�+-S�μ���fFkx���L��8�QW�"b��Y�[7�pM�	�sD�;��@,���+ 8�8`�VxO�K�1�&F�*izĤ�=u�]����%tp�do�������Ð"rLc�K�amM�r\��{�d��-�͎$�2��Hx���O(H�)_*���|Y�w[�'����M�+��@���`E����h�����Ŝ�#p�6I$8k����z� I��xHW���)$�@�TKk�ou�她� :l=>� �9+U�t�\$%GrҞQ>�~M�{�ֳ���484:r ���M����8��푺^�m��ї쟴�(k
t��ضܷ�JW�gp��1���K��nAO�U.��3��{�9b�z%(����
�����b��w(��|�D.\�c��q��8E�h�9�y��Z��H����A힓�����<��d8�4�����5�1j�����Â�U\>���
(�0Z:��;slF?n.�:����~ct�@��}
!�;:�Z�tN�i�om�[|Q3v�<A����5ʡ�*�12��T_�SD{�C��z$��?@�0d$��hrp��1E��f*x���"��p�&h���'q\��	&#��>�A��������U�u]f�|���!���Y�W 4|����A� U�3@�h$*��̌$�G��~�������.	z,��G��ӱ[�����s����{Zt���s{�=O|����h��M��й�+��I0+�K�w-A�un"Q��_�}� I ��
�{8�ͼ�3W��6�B�g�>Sw�$x����(�ի�f|���03A&��}�J֩y���&O �ǁ�0�y�d&��y�)�%S��L^ph�L�QR[�主���ر]8�v~H��~�x&z���9�Ⅼ�����h#Е،F'Q�vb���������g��cR
E����_��5<�@�5����F� ��3�A��Q������|�(��I��.��)�eǠ�UbS[���!�y�� �a˻�>W|6Of)�Ϳe��Z�e�*��E�:Jk�)�x�Ԑ�E�9�!�s�\�C����G�?Ȳ�,�jx�{J�,A!��^�}4 WV��(@\ǽ�<&�3��^VO�X	~�~��'\��#�dt�zr�>��89.Yz�$ZPd�N�v{2���ݚ�����;�+�����Ԥ1 �2�7k���MO(j5��x�i�8��4]�����R��~�63��EKS°e�m��7ﲨ�h��0Np�0��K���9�I�i��8�1��dh�T)^�����K�5��������.��G����8�<�,��ۂF7N�-�#ic7$R:��f?�-����a�`��q��]���:e��1d��2��}�;�+�}��|(r@�.�~zxǺ�'��iȣ8�����EX�-��/�f9�@C�7[�rOR�f�P���u�������s8@�ㆶ��C����H0=�n6�~C�L�?ﯴ/�H~0��q��Q�Z6�D��_��d򭄽n�Z��x$����ZZ��B��鵹���C���XG\SB-�f1F��+�0^�%���ѿL�2���ѥN!5�a��B~���E���2��-�S�"`� ���~*�{X�r�g/SQ���<�ad�}y����D��_�^�!�g#��$^-q�37�-|C#ݬA����Fn��u��1��Rd��5��ڔ
�$���'�r�n�}��8s�� �:Y.q%�Br� ?M����њa.��p���1�'�/��.E��k;?>a3��iW�~�V���#��&m��{���(ء	�I#6��R�ՙ�[B�+�֑jy�g4��\�J�aQ�ЍF'rG�t�
(
�j��S1��y��S#A ���{u�t�>��tŔlh��
��jN��-q��&���:��Cm�^g�=�ۍ
2|ml��w�����&M�>�y�	�A��~:Ŕ�(TW[y�2}sN1fE���OApk0�/����M�6��2���?�xY�uϞ^�"��vA��P�ra��M���*��z���[2����L�sR� �,Q>�`�n��	�_.`�92TxSG�1Yh�X �"Q&�D�;E�(�����1u��@%�$�uS�mЎ�>�ߡ�S2������l�!�-o.��;*�`������;��Di@;���tg=ץR_�K8W�����cG�4�."lW����h��0�n�Z����$�1s8�*W5A.48Uػ�}N�#�1ǩ0��	f��>8^�]#�����ƭ��o�^�11;���2k���,[�R�p_�;-�٣M�y�|�X�/4rkV�}�g퇩�K�Y�w:���h#�0	/�1O��:}~u�^p4��n=�c &��1�,'2�h��sSgr��C���DR5Ŏ#��%�r��U��`e� ��v��rv�}��;WW�ĥ��R�G�n ��M�m��D`?BL9�����o�^�ٿ����C�m^:��ȡt�HGJ͡���_����B���N"��Yg�g��q4~�L��>i�W�_���U��E�S�IAm��Ӈ�E?�u��	;�+2���F�G�)/`~Rnf�'-1��{��s�T�{��w@�0�UB���q�l5�:�����:��Q7�X�L�@V�`����L<7�'N�J���� �ղ�e���,��SL���|�Z�悕�ׂ�R�,��\r���<�)����u;������� ��*�>��҄y8Yy��lƷ���P�S�L�!�ItP62m�@�1x2}%J��.�-Kޫ��v��@:�y��B�Ml�<.o�������2}r��ڢFi���jX;���X�Uk5{f���x�;Qn��)�}��iMM���xv�4�Z�t'�w�\c3��k(�fEО03!�>\����}ym�v��'�7.U�b�&Ɛ8��g�:a]��]�}*�4�'=r5�j�2@)�$T�I�ž��P�*�E��1�$X��J0���*҂:|���v��ai1# }:���'�y.fֺ��QK6r��I~F7�O��Ѵ�<�pQI�Jw�|v��m�8^X�8k�:ڔ|�cv(ҤgRXh'
0��k���Csa�?ے/�)6&3��{x>�Tx�y���1�s��Q�v"U��Kp
<����*�����ƌ%�MF�/��I7֋ck3!~?�[z��/�7����^��ײ:��jE�k��"S�u��I�$Q?�H�A!+;Bv��l���K��hf鿅�c�L��є�GP�fw��;��{<7�J��4;�����%�~�(����]�'O`���k�-�Jn��������È)- @����(�b-�Bj��
zԷ����j��$pk�
&f�ѰNf�H�1;V.�_�T��Ho5�\}dr5+��N?f�ysHPj���s����2��M���dq�@l�m[0@ς�l㓶�r�(�\�ږ9�`h{EY����=q���!	�+C��dz�lj)L7�����,��G��(���`T��gKs�w�"���J��ا�@�#s��Y��'��J�bR�������E�w�_2+������T��8<ڝ�x6=����_:J����@��\ũ�Hྛ���]��}�GA-�(�XldڤɄ5���Q�Y��kv��G  ��=k�"G�$��������H���3Bc��-2��%NO	ɍf�#In�<�@M LR�!*��j0~'���:L�'� ��`��i��(>|�0��C���l�[�0�(f�f��Q�D�������cH,��5������#�rdo�e�U(��'Y\�,<�)\8�@� 7�׉�m�g'�%��k�]�"�uY�Y;YF����A���Â5 ����ڕ�mVhX%d��_%d@d?�?��D${'������j��9���¯��-e�1�~�箕�"�/�|�Ո�؂J�tH�}jg�]x��E�0i6D;�g+��B\>3�
�	�-m��;u4
v�W���ŀ�� ^����~, L�yx`���zN~�� <f�NC����l[�"����_D�LM��.��<�zp�a�oD5V9��� �Bt,A�����8s���-���+��E�If@��F��ö�<N���
P(�N�Q'��/߄�;�bB�8���'mD.`�rC&\�O������W�&�Dv�7n�x�%>����4-b2�^Z@�6��'��e��y�^l.��Zu@ޯٯh��*4M!5ח��#��Z�.����^%X��M\I�DN7�2�ݴ�����շ)�p�B�����h?y_=�����҅c���̓�l�������NNs�� �;�<`Q���vB�rv���¶���4����A���W�#�Q, 2����%	I$V�@�_#���-��	�φ;�야��9�\I� �ѿe"��:��/Â7!�XZ��rJ��ߑ���n._l�X$K������7�}�l Űx�c���|V�E��O��Õ�P�"���pb9��1]�}��`�mn�#�$�Gs0�Z���S/)]��յ�і��8�n���D�T�u��	�o2��AGأ1r���Vb<��yň����ᷯa��`'����h��Y�:��k3S.V!�J�ڎǠs�禺��q��+�,�W�9�*46=;Θ̿6�*�I���c���g3��j�l�6.�oZ�,k5p�U����1x�ғ�K��ϙ���K�R&��X.�	��`��)�ĕ��`yA�xIs�AR��R��9M�q�n�d�j�4�bC0�T�|m�E�-�C�Dx�i
uU= �4��<��ځ�7���F����o����!�r����ik�b��	�����u���^��g!!T��e����Z_a?���@йt<"�Ϟy�����[����u�2��k#&�`@��[�h�{���6��D��6A��`�5�G��:��1l7�x�(�֫-�V�J�6�����2���S軛�;w�߀�i�G(��h���V��cK9��ҙv�8,٩Uݻ/�$pތ.[��e�e��@[Z��u���W��-P���-��<�	�l��BR��VO�ꉉ�7���"�,��r��J�E��9�}���I.�H]Рǭ}
�jk)P�2z��|�ӳt��t�����p��ჺ�WE��p����̿���.�8��g=/�š
��=�4"���M�)qMY8��Dr���ՎZQթ�fs��A�+�y��Y��/�ҁ���|^������5�A�.F�o��䜿C���� Ю"h�bB]�L��kZ�oZћ�y���>��O9[N��>+$Ҍp��l�7s�"��	��D��kB�'��$�S��sR����W���ĩkv�A0aZ���&�����1>�@ñ�����	���=/_.,�2��7�~ul��H�m3�x�B�%�y�q( �Q�]���q�� ���8�����]�ܒ�m^0Bv!������&���:�@*�!o�sM��4��Սj�]��sH0lBǹn:���#fx)tsf�Ks��G�#>�̣�}���7o�:G���3��4c�2�;�%ՠ��%�=i�~�Gw̓��YBVf��̦4�9�}7��e�ש�<Ag�pc�A
5_L+��oXA�,?'�Q��b���o_��~������!���M�eT�������ܚ4 
����@g��u�#���&後�;�HJ}�tM����M��R^xk%K����l<�Z��kѴ.Ԕ�@'��H8�%�X�*�v��JpeW��~�N<�Yq�$i3XR�w{�V����Є�(���-��I�I���⻚o�[�%�sl����Iu��zv����2
,d�\��1�!��R\�Y�,˜�?�bU�!Zp�AN��y:|�����RsJ��EMxp�>�mq ~�]B�v>_3�N�j!�U(��I��#asGv�/#"�Vk�:Mi)ye�͊�=�GX���H�'}�E��h�s_�g�x��.4Ih0.`��*�6�P!�}�lU(��%�kF�'��MKu����r�O�>��	�롾�ȶS���F;�pc
��|�n�v��YFc����B�mI��h���f�kz�{�{9�	YE.��JnB)��	V���F���l?��E>}��;��I�Ǝ�4J|��p	A�����1�H
 ��"���d�ޜq~̌�	^.V�]J�o��Z
���{��'�#	!�v�GZ3��*Ȟ��w��,A�;�7M 34�
zo���U;'t�)���?�J:j;o�)n�Q�#�?���"����U>�:�3,g�ly��ޓ k�?-���8	��JV�\��H��c�#V�?��M�4�R(l`�z��n�* =�5,j�Q�������U^�Cűl���}Z�K{q��r�a~�.�*�B�'f"����
���*!��r��'IP����R9��)/�?@�2G��o�O%Q�f8���DM�	�T��ߞ�h�Z�ɂ#t������/�ta����2v�@��_Pcz����@��k'ue)R�յ�����p~�`�w\ @6/A��00��^��A��.!Ij^�m@᠘�"�6�%�'��ϗ���EAV�#�$�����;�������Aj���H���P��l$�J���֝'��7��J���%�ݹ@��g��}��.]��7�KZ%+K�lH��a��唅��e��)ϵFvF��4R��3<mT4�qͿ<P�����
�M��j��*9�o_K��6G�'��cQ6�M�mޢ5sh+�N*��=ܦt�2@�,I�$����g�>��7=�x�͘�x�>O��&� r��ȨySL�xR�ѡ ���͗��G��DGXQ����Xs����hF\���"z� ͔KT��y��v���&꯲������w��7q��Q��͸�,��=,�Q�2��5����p���)F*�`7�^���Q#�N����zB���E-(me	��&�č�A��7����,u�_^�?�um�G���v�����G%�߿�������$���S���]Lآ]���t��'��tY��_��s\#����8!�����+���A�G��pƱK`V��9'/2m�^�m�0Ul�hB*�0�Hq=pq]��x�2�r�����T�)kRUSd��F|��n�e�o� �z�W��n��]�7{�_I����/߆fo��D�� ��V^�
'�#K��E���~�i�?���2,*��ʀ���i�*]qI�K=p���#n�5������obj�bxL��>��9Y�6*�����u��!���9�-�VS�g�RE�]φ��+��_���
0=3�b��V]�(�&���̍��As�:5?�R���Ӽ��Ōh�����%7�<�V�����*�<ML��k�mC��4�[l7���{cZ�c������3�&��hv��x���;��X͙��z���D��ȆO�`�I�$�t�OXB�&��t�yp�ǣ�|aP7�7�}�^��R9��lO��"�HRZq��,s��㈯Z�&&���	i'�:Q��x�A�`Ci���6R�}�6pF[�zLe���c.9�:m�'w+ou~.����=L�LM`L��֫E�)K�?�/*�K�Vߛ�"�_6��{p��G�\���.O(&���j�b� m�z�]	6��F�y\W}�^����.hBӚ+��K$@��	Ɏ��{l�?�F�o9���Ӵ�%�������_�N��*�-�.(�gc���Tkv�o�J.����^��W.��B���
�3��my.h�$�F�X���?��r!�| rk�5���%��c�תE�U����_곃2��f?�h�&@��颁��%�[)�0�3a2�g�nGf���!���:4~{���l�\L�㨐���v����j~�)��C�Z���L��E�ƍ˃��L�QH=���D9��yk��<9�r¢���ɯ��9������ J��J�)|w�ҟ�\����]��~��2Rm}�Bē��,��
u	�uPL�e���B�:$�x�l��w�"iͮ���>:�vc�^�T�Tl1C�"$^�t����n9���6������>��Q�_�o/�"���V��l&��NcR�f�#?��+-��
�q;�n)�axvs��L[Th��1>t?&%�P���
A�e������G���4��-#f�j}��&���m���I�\�L,N)&F����S�Q3��99Ѥ^�`��@5l��8�R���;�w@���3��OVb�7ޜ`�Ä����4FB���Cb�D���%A;F���Ę.k1�P�Ul�O'�(�f.d������F̏t��2v���J�,y3�H8K���G���,#�4:,<Rj�?zNr��P����`RE?n-�Q:�r����0P��P�X������\���S���św��8V]���J�"MP���rD��M�3	}�In2u��������jC�O�V[�ޥ���bUc���{���͍'�-�7Ů��-X��L[�0�j?a�jpNzM��E"��ҬÝ�1�k��т��2J����o9�^2���Gbl�xc����M��5��˦Z�Y}��U��`2��b���L�1b�&
����@�^�Z���' ��.S�ڂ��]���mȡA�	�r���v
ok��tOD�A"N<s�A	E�(MS?���PJl ��}˸�|��L�.?�&�A��ǉ��h�4hey�-�=����R���0��D,�7�o��i�{v=�k��129�1Ɵ����D�`u9z,�՚L:�{''`*G�6���Hѯ��p	/&��� ��%���g�Lw���I�|>�3%��]�U�b��/Vl#0�<݁e���a��|�U�!q�-�:�
O< �,��_�d���Y`Y2��6���C�y�J��(M��m&�JlҢb�gU�-WN�v�s��$|�O�eD[�2!��J��`�_����=��;݅�9Lu�����zȁࡌ�7˲����l88S"�>7ğ�<6��ab�0.9�jl�لᣕ�&�� ������m�`�1x6�뷋�xA����(����
������}*�P.�����)�aA�,7�!h�vi\`��UI�V%�8�������+���f�
���:1c�n�����
�;��n�<�˝�z?�H��x콌�eK��J�R0g^7����4���#��u9[N��?pp�>�@�i���ҕ�K�l�j�#ыɠ��<2��#�a���1tw6�$J���$�#�8�H�.���]����{�	������"[��"�[�:t�WUh��nr���o���1��ˎ��)_�#������� �g���׍��np$�V;��]֡�������@]8��{"�䓌�V��i�r��')l�\%�j{��l�<�L�D�7���r m�1��c		0��� �g���(�Mc$�T�4�zBl�p��yb
��m]&����ej�����`8\HkDy��^�z�<fe۫���I�
[��a��/RЭ�����:��Ý���T���Ȋ(1�}����9 ǊU	�~J��#z�r�:'��R���g(i�̍��MȾjTJr?�D���2�d��Z�!��z��Əh� �V�LT,���~B�,r:GO�N�v�ڳCp�n����F�a|G�'�+6_[�T֦����b��y$��5t�=�Il���AQ?@b�D�on5/�>��<g��]+y�����m#�-k��y�z���pVX�T`Йh��/����1�Ӝ
���)���x͸p�����K��
�v���Ht�~k&��˾�����t~-�����p3�r�k��V����2�	nN�f��ei�\ūm�J�^�!9o�k���"���1�����q�_U3Nf�<�Oڝ�T=��>����ݜ V�'��Z٭$נ]�*��5�,2��b��	͘�&T�6;��  �v�*$Ė\Yxʰ;�chD�d=A�1�(g�ΓcA�؞�#
�3k*�1���w���@v����+�2  +�4ج�k���@����]�#@��	��Lg���yL�lT^r��.��hv�.����f!C��ߊ�]XU�hj����с7b������>��0�\S "_��&Eʴ�py�Is]^����LF�4���B���gn�XS�h���=���'��D���2";���M	�?=N�wO�>��z%/���	�;B�����0@I^H^cڧH@o�C���?��d@�B�ҞX�;,�^g8�A~�8�dz�~M�(�CD�E��r$�>�4�I�/�m�Q�,f��-`�p�N��פk�
�fȣA�7(8�A��W����	��Jj�狚1Rm/I�ΰDKtCx�V]��+�.N�;�m��3ą-�=��ҩ#�M�+|�h�۫��0ut���hT��:�;��_�(�W9��"iu>ps�)8I�笯qf����X�A�2%�3�挒F�׋5dP$,4G?dh�4�t�^~Z�;^��>����-3�#Ό��C! �K��d�!!ݚI�ʽ���H���8o�����KP��t�g��ݲc;�H�Ϻ����j��)�!�&��� U�	��$WB�FJ����e�^ӪE�3U��%@�0d�i8<~c�W?MA�#
��L�!��l�I���}Tb�-����B��zyitE�3&��c�lπ��m3w�Cri���z�,qȨ�h�W�t�6�P&T`�Z��H�(d�\V�Й��:3�Tg,�fzG�**�Ӯ"�j�8���o��~ �c�z�~2�$A1�~�u��_G��|H��=���z��c�Z���Ƙ��1�-�,��ó��j6���N��"G�a�(��Q��a�y�����v��f�ߤ����{�ڣ�}ەi��F��!�~��8�[T��������k7�9�	����V&\�H�8�@T�2�����!����R�D��p"�Hʿ)��|!t����"����N�>|2mj_���o)��wùٚ��XD_��o��Pz�u�i�~�U(\�?f�0(�RV�.����w�:��Ӱ�FĨ��Q��8.�W�us�4��b�%��bq�*��F�*���d-�@�}��e9�A�A�0�5�Ħ��F���BhX�n=��$ީp6�9w!w�J��OF��]����E���Y:��sh/�_��*R�M�)S"s,�W�?���?CߟN?���A�6U���Q���Vyv4��)O�Q{��w�E^�f���޺�>[�n �W��ڱ�T_��0�l�Sn]��N��djXʸB��J˗���}W�������K�d��T�d����)r�B�h��~t����طL	�Y�>֝�KW����le;xң�dqo���k�xB�-\�]��ԏ#��ғv�����b�ѹ1�Q@Hg]0��򌧴�Q�L�Ү �e%u�hl	����{�ǧwd�y�Q��w@�U���	!;+�~�'V�W���cV8���O> ohP~�$��ۑ�4J��̦��=�������˺���vf?L��%�`0$�n�5�^Ã(P}��RM�T\��ݬ�O��9 	�h�*G�X G�L��6��2�Z��{�J]۸d*i�;�яW�,5h�3k$�zS`�X�b̄j�n-&0Q�S%�N&ܷ��+����+|UR~��.[�x�Ne�k��oFv�������X�L;q`ک�=�wm�|�Ⱦ�[#�p/�!C,��:��՞�;ԙi������NU�g[��~��^v�#�������d  �𧶏���w�,��1�I��b(	�Z��o��1����p�hrsA$��f��3�G������?���K�4�i?��G�� p��B����5�f���W6�s7ۋ�l�(a@�t
K�z�����q�b����H,��B�vԸr.)�7w�/��oƊ��I�<�e\�˱5a<�?�k{���F�� D�%RC�lgr�6��jj7 =5H�����g�O�7�P ��S���R*�o�W����ɣQk�q��oҬ=L3D��P}|R��A>�)�%�c���������ߚ)(3�JF�G(W����?���i^�Ic�����b��@������L:9�3�˃(%�[Ht����r��q8fm�~r؃c,��C�)4\�����V���ؙ(�;�~ۊNx�ʿ��6z���k��W���{-�@��(�����VB�+���+�09�g�{2�h^K�j����~x���ɕ�u�hz�m�����B�/}��v��<~T�2�5��#4J7�]������L��&CUMiVA ��9�\^��ݧ4m�>�D��_IvuN���[}Apu<����p��[ɟn�W����Qbg@icD����J@hP����M�h �-H ˾M��B�cã�@��ۉ�`;j���m�jV~+?�OC�?
9�^>c	�oL�� =�Q���;gڑ�Y�B>ܥwfD�d������"���f\[����;�U�t�I&�Ė�%j��3�O��{�h�*�z��e~+#H�J��f��T�I�p*���/���y��)@�9�'S/Z�E9�v�NEq�%+멉b�SE��-0x���D C��B�{���A�߉��:�{�1H�邫�b~�ր]>8�]c31�!HI�8��E]��LIns ��B"����$�|���Fߊ3��[%��`�Ϭ��uU�ǳ�f�$ЌK�1��c�{�#:�0HL V���m��_�]���^��ɲ��R�:~�<����Fb*�usp�_lb�cա��8t�$dx��+XN��AG����2;��g��dyD�w�qť���c:wQ|X� �{*���=���5�b�����̒NO�2��a`���S�"Ϻ�{�@����h��5&�����Ѝ���yG��P�����>�Y*eii�D��:c�������6H�d���=ͯ1��Z����{�U���I�����w��"�~��Z����J~��Mܬ+��D����x�E�-��$�����uՄ.ޯ��
�O��F�B��v"z��y;�����yj��Y+��dF��-d�E�5�-��-C�=��\��;�к)���`�M]uk��s+�豑��g4�ѱ	�9<KJ@M�Q������O���wA�'!Z=V������y�K1	���=tn����������ݷYGڨo>���n�ָ�V�MƖ��L���>H$�������X���>j�;����Z�I; |��bA`릕�odS����!���TtB�}@�E�����=�Փ �ee��6f>�������U@��Q �j�[ҧO%� +yk�O�����p&�,�%���L�]�\�	&w䓗��ƖnM<�<H��y���`��m�i@�Wޅm�.��5��3vI����˭n�P��A>�Ұ+1�Go�C�A�%M����Z>.��<��ŀ.��c-��wik�m�V���o��X���,C�v^���i�i"��eٝUfv?�t��ٌ�5���V��B��$�Ǐ��h��� �«�^?>���UȄ%g!�~)r>�Ye�^
��Ϫ���O�b+E�y��p�c(9�Se:J�>j)�?���o��e^��.�9���6�S�A;�<�s�{�r�xO��x~���(�R��0�.qk�㙻�.�c���?g���� ����3��P)����;��[^�,BpB��܄h���}���2P`�P��K.(NG^ �~ ����u�o�k��^C��A�0�ʯ9d7��:kke�t�@��m�d
b3+bܲ�'��)/�^\z�Q��-6�|��L��yԧ'�m����7��L��b3�&�h�U�������Ï�\s8�����ެ$o�XՋ����^~fz���·01�/�kS�{�ܻS���%AH;���=����H�ҿ� S���'Vp\��<n��V'�TğQ���lnfL��t$�����#��������t��vv��x��-�̈����TeUb<s�~^Y�D�N�W���XW��	@���}߻H��'�.�� ��-�`�@��{����-A9�󭺟��I���=�����sc-�* �'ܱӧl��5�w���?��7@0}O���l�l�X/��. ���W�_0�s��-L,8��U�+t����"����RO}�C�$g���.I≞�z���>xV���a:����Oa*�g�R��W�k�X �Q�� ��^��N�����N�\����E��(G`���������Q��y�]���f"��������GGuʠ䘱/;��#1��ݏ��^�|��zz�[7�x�n/m���8�h|r�,\?FC,�S��;����Ԣf���*.{�_ƭ�'?���)Ep�z� �s:}H��ӣ"����uG���E� �8`�����D����HG���m���N�.�D,&��C�_�`���T�K:|c�$p��D�|ܑ�Hs���&��Σg��'w���J��H�=B6Ld�ū`G��^Y��#���#�}�� ���We��`]��Ev�Y���1l�n�Ӯ���=�L�u�0�[/ˋU�~�:àF���y����Ie"�ri�%G��6�g�P2h��t�W.���?�����қ����Bӕ;z#�+W!ͥJz�IeL��y��Z��9<����m��������Ʊ�DԪ��Ĥ��жy��x�c��z���X��覅J_a��6@�K7�8 8��t�tdK ����aD��&pG9z��I���F0�t,E轢��|�"�`�1�	/_(,��;S�n�ˉ�$�^�6ړ[6�j�O�jV��2�K��j5�dm80��{ɻ���l��齔:q�|���%
�\9�eD�)(��Ƿ�9a���.��rs��瓎��2�ӆ�jο����v�x�P*��� �l�Rf�>�����ۤ��PeME�m�=yb��v�TqG��:��FZVO�C|���£^�ͦ@$��M���B6��?J9�zj"~H	Zh�H���;2�K����O��l�gL�N�q����CH�sPg7��-٣�`>�ę����Ⴅ�p��ni��ց}xse~�Ǒ�x�0�Gm��-Y����0F�h3y�ٌ* �o*]̴ʉ+�X�V��ܧ�0��e�jB}W����ǵ4��OK�̻��<!zT���W��Y"�h�%�̯���(���X܎*'w��EL�n�5D�0'6���os���G����z�!�}#�^����@z���FJ{�α���[@OE�eS���9�wn{J3��U:��������Py�����K�}��B�9��q$�˩D/oؖ��8F�.&��3��8�3]�-J�!xuwM s=UU�DyI��j�})��B�꟤g��{NA�s�ecl'a)���b8$k$�"�!}�px����h�"n��A��9�d���\�����/��L�/L��|�?roh�b���+'������
x�9��11�ϩ���Ϸ�94Њ���9A:uaE�
HS��Z��J��x��9F}�4ו���w���-�l�l�)G59aK=1Ψ1�1�nF+s8���k; �Ot�ί��\�����X҅��o�bo��6y�M`z�*x���	�LF�_�C=Ĝ*s2=2�|��|B0�UA��J}'��w
"��?�?o-�1}�>�\�NJ��;.MQ�\~{�IJK0rl�
Y��Ce�����;۶�m�N�.(H���n��g¥e�׭`������ИZ�`�+��@���k����\ϧ�Fkɉ(�]q����-�jtyN}v=6t��<�	���`o*F���%��Ձ�R��X�d��yD_������� y�f�"����mbbmG6*�4�E��7Lg�n�Sq� ��Lr��N\�*�|��b��d
n�c�r�܈��֬������ю�G�p6dY�eg|ǲ�]�z7P֋�Mj�Gi�=	F� gH*�?�Y�g+����g�'�{�m�I�Y�h�l'y{�~8iP�]�rj����+�3I$���q�-�L_���"(�҅ai\d=�w$t�Nߓ8\l��V�Ð��H�Lw^����������)��ϗ���s��u�g�d�M��$��e��j�r���N4G� �$:��s�wd_<��<��Ԍ}��D�%i����c��D�J��3�I�]Ny�Ș���8zO���p&����E �|�3�����֍;���e�t/dܺ�i7�W�S>X	���bK����� �z�Ӝ��六��DP|ġs���u���mX�����9]��>fۯ�t2�p�:��/������i~c4	�j��O�v8�R ��W�/�1��ϖ�5j���d�$>��	k�B�W��i��Ϸ�6��'Kwx��p�7E�����N��Q^�_��i/�\hd�J�f��� �DS�S ��_��8ISL��,ְ��:#��-��+���b��*B	��2��M&Η"�"r�1����?."��֞S��?*����������	�F9׺RRA�ƺ�ϰ(�'Iu�QH�ϵ�m�Ug��a*�<�|�jI�%[4��ul=�<*bc�.��V��!<�(�
)*q�T~K�"N�#���~N��)f���L.��~�A��c炶]B�T6�������x��B�����G��##
Ǘ���R����:r��\��`��G�2Izgp�O�'�C�fc�%FX�F4���3=Q�I�1�P��<�%�\+�@���\���R����,�Y���̟�y��T�̏���҄�T��#�K�~yH��A�ۂ�'N(/��l�gW��?SL��p��ީ���%����B)Q"�dv�瞣�bo�/I���g�E�4��^�Mt7o=�ug��Kj����N(�R/--H���Xp_C��;�j�͋3V}౗��+�!!��ͷ9�=�0�"����a9b��7[&':�bR�s�9��eI4"[�4�[��Sx���:b�N�/4��Q�]G�"��,����
7T�0<9�.�hT�*#gt�X>� (�`�ͥ��̸�@^}���1��b���`;�@��FI�����r���i�'�%f�x��K�����}��CTN�V�?Ƹ�����W�j؇�]5�����g]���8��;R{Uγ�ׂڲ�[G��LT��p��ۗc-� ��>�t�y�����y��P?K��|^d3�ϓ?滁�d�[_�e9&��0��T��Er�h��=�g��^�45VTI�5O�:�ɂ���:C��.NZ�f0��Bo8�|5���,��ҹ'�ܻp�]�_YRJ_�&Xx*�� ho��	�w��d��@�#�D2�����Mo)�fq�Hs������
����Q�+qZ,η����=�����Fy^��Ǭ3�G��`���gr�v��G��� ���aX/�.�����]�Tbk� x���	�y%}����K�@9|���\9��)��\fbE[/��JH���1�����` ,n�?	� >�k�	sY����熾����V��m�y�SJ��#p ��X���g�,9
�p<;�h�b�^��Y����Omw�x���gM";)PB��C��M��Q	U�A����(�>t$����&H�D���ͽ����r͈K�>�����&{��O�/+��0�㪁�ɼ������J,eVc�u{�)�����쎩�
���ȠX�;��_-!�u��������z-��͓�SI��y���O�܀u��fJ�*��&���藍8o�g���P��������&��2?aA�=��\�XU� =$�W|���x��h8T!��� �M����x��a�8u���7\��[n�=�OXGl��2����\R:���E�7������˹�O��Y��� ��ܺ)~f,yx�>���1x��׺�M1V���g��`Q��Y�J��9��gz��z�M�����؝6�k�^�5�Mm�����AZ�8/Id�r�a�U�3���l���x�c�N��w(�l���e2D5>��#�\Ѥ�즋���J��5��)2��-�U{y�D�LZa��|��_�(_����7ܞ��Ww��N9²�{Ý_��h�,$�}u� دXS�q�^Ѧ� ��<�UeACi��.�{ED�l�	�.g��1�&7=N��qv]O����Z.��1�_�W8Y�p��xa,�ɏ��l�9�clvXF�u!O�c���I8�����ٖ����6����}�b���k`Zs�EOAK�"�y��h��J�mL}jC�x��&X�L�۹SZіR�s��8{��X�//�a�S-�Yi}x�&cQ�� D6Ζ\Uf������.@c���a3�,��
E�?
+v�/H��&����v �W�('M���(k�fm$�vY=v��;<0F|y�?+bL�-b�5�
��K�" S�]��v�6+��\zu����� ��q�)�+��j��3����D��ĈLH��?�q"����#㸾�j���E��"���K:ؽ�)�e��&K�ڸ-Jjz�q8B���h�gYf�5uy��+���P��X�>,Rnxi$�la.dڈ8}�
�c�;s��*%.o>������J�����)�3���^����R!�W3��p���i�����+^� Ïfb5��$��(n5[�ο0���>�zޠ��ݮ9�5��y(�c �'��6���o5�F���72:4�����^yE�M�T��>��t�]�tO|���<C����\)�-�Y��;ȷ<kNmϒ�`�7/�b z��V�D��������ֻUp~�B���$�0���4W T�#���M)�ꈰn�B�U��P+�zy�/y�f�b�6����Ƴ{t��W�)�w˃C����Cv7���U=��a��)��-j��˰��� �\�P�e6�>R7��M���x�I;D���]���5�H�����Ҍ��VA���O�Ңr���6��[KLv5�)d6��\t�ޥ�aS���F�@�����H��B��&÷�4�M�A2�s��(>�<�H_b�X�,|J�����u�޲�X|���wH��0�_�yn����g�2	]}�8��R���GZme&�� ���*/�{���/����q����К��^ʃS�,ϡ�l�����ei������~K/�f��R�c\o��ڛ]��x�-����ю��²Ӄ
�M��O*[&��Y�荬����֍�tI����u��=�@��!�+E���)�*iY���~CqcB�Q�k���\ߣ�[��lr�Ȭ��]V���� 2����� ,t���Q$�YVl����B �K�~u���:|��\#@�T=���t-weuK娶j9b tߩ���Xn�/�m�&�al�����u��'�%ͱ8��>����{��x%�{�,�}CH�F]%�ױ�X��aٽ�0٨��]�̸G���'.��W�)�|E33]#���۬��Lk [�)�h΅�*�CV�Ƿ��k� ڏ�"|ߔ��V��//���.f�1�q��Y҈Dg�A��ռh�4[�����H"���]��ff"S����P�B�.
ʛ����{�3'��썆O!�(�^�n�)K)���9ի�P>����㈫��2$��ՠA2�!{����n����pl~,T,=~}g�v�˗��:e��@�4H�l���%�?Rh(Y0��<��%s o��G�4Fy�SޤzJl���E��/F;(�i-Q�b4�+�שH�XG��v�L&$+m���Hmd�[��c��Ռ !u�K�~��0�B��M���Y�v��b󞪾�����|mB��]�<���@�Q��
*�=����� ��k�w!�3D���I�u�SF��o�d�#BˉK�#睙�5�d���1'���>y?�|e��6`n��Q���Om���E�k����w�2K�-OG�Rê�TYvz���C�!&=����ó����d�U[�Ҝ��w���Q\�`Dd_�8�9����$���*����S�/x{|�
�����wFp8;��l����@?���k���m�`��w��9�\Ρ\U��Ƃt���I�`�u�B��G���O�GeP�����U���E�TS������g�z򩒽�Y���C�"�P��(�G��O��:�Tvݗ�2�v�|�����
�9���kh�R�M7�W��طw��ٹ7/(��;��ې��d������a�k��c�����*.�F�Y�`փ�k9n�T��[����@�J��Zi}���v�0�N�G<�V����hI�Ud���R� rU
g]���'۝A����2;e�U��w|!4�׵,M:�����x���.�KV��_0Ƶ�e͖A9�4����ëͳ����K��BP�9fG�y�.���m�c�@-�v%��2����Q'��w6A�М)�/๭	2:W P�3! n�Y[�{�A�G�n'���zW��h0�*�⸅3ꐾ��視`7��]�&���fU��L�MFy0���p�:�<r����Iv��`Y�$������_r$I��W �E�+�5h��ξ�u��b18���IC�M~�)��$^��h¹�Ƭw_��~�6ǩ�Rͺ��#�ӻl�N�>|�<��	܈�3����Ԟb�qx�ò��	�n�uB���#�^Գ�\ؚ+),�N�\���#k"�+�dS��q�z* �q����?4���fu/Z敖l\�.j�$1X��e����ޝ��<��Ƒ �x���b�����\Я)<k���(6v�YamC��m�韑zd�jO��}H��A�Ge�5��%)���6�UI�^�2M	�P���{�):|Gmh����	�<����H;h�0/$Oލ�$1���������uǓ8�0ޫ�b\���iA&b���4����@�a�D����d_�ׂ�S��V�8ƾAx���1��0ϸ�K��y�P�(����@tg�Ĉ��	�h7�	|�]N6q��lRlɜVNܫ�a��d��7��["FIxZ��Ű��#É�t� ��6S�B	ҷ��a��t����ko�H���ɘ#���A!ɯ���{�0W��2���%]�s�h�Q@�P���Zo$�3�}��)��?ȟ~7}=�P�1�Y��V8+~�����:�)�WD�X�j���7#W?��_�R�dy����n�3�x�0�����o��X�2J�T+SiP��ڱ�= �r
1߬�Yw����r�`��~��V3��kA$��3�E;�,/�]�	�YP�]� ��Ă_�UAi��E�[�N��M�xꁃ|̎yvQ��_f��g	�ԵM�Q����8/�����B� wǼɗ�����Tm�+DHz����[��g9A����a\��m�5^�0ǫ$Ђ[�a�H$����*DQ�R�Ѱ<Zώ�^�qX̙�o0-�4����6+��#��}p��Н��� 4���ZW�.��`&g��x�T��JC��H�ؾ�% 0Mt�~oNq��t�Ɍ���2#��*r)���Rv�c�&��	�l�!��xE��s�_�^�]m��כ�Z"Q�eʉ�!{�_c�rf�ÒWҁGX��$=���j-Z���<�_�͚���M��������=M�.��;C"N9�^����q2�o��EE�a�#�	��Y+Vp"��-	�m���JK���I�L���2 �X��"#t�)>�Q��޻|�[�C�I5��eN&&���9PK�#�������l�th ӻ�Ҙ�ӎr��'��xZs*�pv:T��ov���~&!�ZO�/pm��x���k3�%/NA��M�*Y���)�P�%d�FrTT30	!W�}|�����Z��/6�V{|�/��w� \����������[7	r����b�[髄�� �m���ʷ�8k��Uȭ��B�o�~�"[g�0劖�e���V�d�~3�l�P"��o	��2TR>�0���L觐gϑ�W��Zh���a<Fȅ.�09JD^ +X�2 Ҩj���ꞽ˩Bgٹ�if�z %��C�|�ry��ݐ�	�Ǘx2*R�\��ƒ�U˴H��n��]y|�<�c,x�I�M�b��7�D$�,�s3F�� ��6�y�류�ej,:��"�EK	���cL
��I�x���TCY'5�b/�;R�t6�yxU�>��:TZ��t�8r
FM��%:��z�GP��ƛS�-���>?���3��ߪS�G�����]�q�" A����(���)�r~�	��RG�&�!kF0�D�4�/�J��8�K�{�/⨸J%qh�d%�l?������;�K���&R�G�՚��ٹ���M�0����j�f���.5wV�\����=ˍE�T�D�y�n��g��D)���S\u��M?YAx��+�XgQy�I��D�ս{��ٚ�s�cVY녜��Q@,����H��``QS3��7���z��Ә�F-ˠ�^��p�>�6�T�Y�T�4�6@���S�e&���;�,��g͚]APrV� N�u�(Z�����mu���t�4��!LK����s��T+��U]/5BH�V3�mK-ǀNڍڋ��iP?�ּ3!�����E�����j9ǘ���±.�]�/��	Qo�`�x��2�@X�����
�r��g��T��1濕��p��.��' .��-uo/�czIh��Xuû�u������(P6�������Z�;�&c��P���O+�ټy!]��N�ub��v�Rz��i�H�s]�S�=�.q�Qr��`iωQ?�D������@<���d�nR"ll����\�Yg�|6�݆��3�<�O�� �er��5'��q�i��YU2�qw0W�ޗpu�3ƶ�:�q��1��J��<�ܠ~�����^.7��4�H"�<!�(|	Ȝ��v���){�&+��o�|�\i�4h�Q��`n�c?�e]8W��ɇp���yiE�����O�G��H���M5����qeC���<	��ϩ��[!N{�){�2�g�(4W��>�u��b�͛$'�q )#���J�Jk�M�r��7���f&�-jK=�0I[.��#�t���{�?ٽ*b2*�S�������zMScp[ 2l�l����������qczY9�g�R���Wf�Y�a���Xy�`Q�{D�{�:���D��}�!f�Y+�c�F<QKv�t�C\I�A���At������w?c��Hw���n\��U���i����7�c�N	W�j{*\�=��CAeO���v��j�`a.��c�f�P�p?\�y1�{���ͩ�,3����
�������_�Z-ȥ�ͬ&�FT-||��#�<���S��t�
��y,��c�ouv�awm�=����������g�s�&�^�z�V��a}�Q�@/�ȫ��ii�?�ɰ�1�f�OǷ	v]f���.��{��s�! K�WKS�:��5`���r�9a�o$�6l|�C��*i�<ÜDt�i��/�k�+ث�O���p��+�����]ж��$����B���>@�nr��T�G=�!ɷƜj�r@�fNEz
��s�zb�]�{0�2~ظ��@Sš�c�m�"��;�2���+���'�+č7�-���k��+5$�n<W���Lu�
�A�tf����:{\�)���G>�?֒�M���r2^*5���:���M��PM����|L��l'���!kD�o0Q��͞�l�nR�e ��3�
�\>��,W�س�����*�,�#�S��(eH�0"eP��&u������sv*��=��Z�37<�;|7��Hq�[��������.��3�Hc�W��<���S�`PT�:��Y�"L��1F�'�-�' ���u�\g��o�D�߹����o��9cac(�����]��Qke*�B���7u3�O�x	��po��x��H�q|�Zw�C��/������67��!̚`��R|-���lK�Vcx��h���<l�~�B�:j7��z�۹�/�`Tώ�1��&�j7+�U�{{�y�����|�3�mb�����-���0��dU��f�����}���fC����"��w��˫�%4f���
lf��ⴏ��^��sO.�p�9�&=q�L��Zy���(x|�"M���y�ITԞ0k�?ܿ��<&��̠��||�v�U���wj�3�t#�+8��T3���HS����V~k,\�̇��7m��Y���݀���A�`���@�����[����uu����=ՙ�
xڐǓӯ�3��ϣ��� K�AT�!:JU�cI5�MD���MY��Z�2K�g݅LF���C���q�ba駴�ʠP���ù-�c�I&�jNd��N̶6LUF6��3Rlm���jZ|ٱ���3�f˕U9�,W��D���2�I�d��r�/�n��CU�/b�hͷ.�ܥ�I\�0�ǣ\Wta2��yW5��n�]j"Z�dTH}��Z1���).��s��&�p��/qu�Y/��h�u��;���BB�?��3�g�j�Tt�ZS�S���6�88w�a<�8�97$��]9f���-M��� ������RCR���-����f�\Q"P{$=�4���pF߱�Z�W	����s�S��Qмx���i)1��N�B�j���&����� 1.��ba��|AxQG	S7�U��1�͠=��-\�i�,ªЪ��~~%��~^� \5�a��圵�-�p	h��Q�"�jؿ>�u6�G�Մ#�?��;�0[k����3a��a���}��/ypB̺����lŔ�:anNR�'��׈�g��/EĪHm�������D�@!��0d1��)���|�Y*�pd�ty��l7Wl��ݏ-��N������$��sՐ�\��PMP\��^?��_c:n�vK�`%�-�A<�R,&|����pt���/��;*m�o����]��i�@|���0PDqE��__� �G�WMp�k[��P�0���wύ��Z�E�,�B'I����:DE�i��O����j �5�^FCE贞Ƙ�.�E\�y�Xן�)�u��w2�Ǣ����p��4Ț�e��E�wϬ�	p"n5Im��>�4y�����I���q�b�,�E��j��ܺ�9ϻ�ۋ��r�M�Q����ݳĴ�@S�Cd�C��RP*��G|_Ne_B��7X_S�cS�~�&!�"��M�~��@UY!��,~~Β�T;z�S�'��~IE������P���0�ܺ�Ku����<g�q�R�@���I���1w^�̀܆��_��b�N��9`���2}�]�x���z�	r���&��~�d����/d3b&��P)�rY���S���%<�zTLez����M�J� ѓ"_�Bڍ̺�z��=a�1zݤ#�����xMp�q!F�D���9� b�xӽmm��c�P�:|�?���dO�ǰV�Q����f(]8CIi�Oq(��b)K��@��V�4��X)�r� ���J��1ժ1�w�wnZ~��Y�1�Z?�F����p��T������}��@hl��My��
=�"�z�Nm�.���4F�qo����K�肁KX�wO�@�2��M���g�.E���s�Iw2
���]%��(c�o�Iy���]G��M�C1�X��0���A4/F�e���
��!��\��@p	둳g�*~r_Ĺ�SOϙ�@�}o�G�_�*H|X�]��̜_͕�H��Yt��"9�1��<�hZ����-�Ʒ'�jk����Wʿ���\���2�]���UPV�Nr��p�ein�Tf�V\�(n�R�Z�l�?�̀���z16	<M�~�Գ���&�iA�V���?*�/ 8Π����0�r��z񃞘��Y�o]3���.�g�!��P}L�C��6��r�}�{ m���mA���y(�Qn%.U5ا4�;��ju,H�%bq%,��)���qb$�v��-��_��"'Ȩt})��3;�/�,?����������~~�q+�B皊�	��vO��F�3'�e(פ<t��甇�F�)0J�4��r�1W��!���d"տ@�a����4^��C��$��b���L5��>�㒷��3Q� ���/J�?A\S���k���ES�g��HnP��iCLU���kw
v�����H����3=�CQ��;C[Q�(/#2((��v���m.�&.��`r8�%��$A�b C�A��A��s ��o��i?�ؠ��?*���L[�i����+\-	���E�����A#��Q�r�0�P�����cO�]���k:Ȣ��K�� v�g�<�S�~d_Xa����:B��v���m$�$��h�)p����
"ڛ�0f���ur��'Z��>�ү)�c��c�j9��&�\�'e�\��aݼB:��[t!r��y%��s�`A�	�jZi@��:9�t�����(�n�����I+t��*z*&�5�秱�xzE�CY��{��٘�N�Ն���8{HB�A�N�4O��n��^h�b���3���������&1��;�2L7�N]�q�OO�ь��5/�:~46�lM�! ��+~��-�$�)j]��36�=Ư�hE�κ4ϡ�V����;Ia�2���̟��+A���q���O]W�ı�d_��V�]���][2�l`mj�B[�v�)���y�\�i�k΀6��b��n�(A
?�"/	2j�W+���Y��U��>���g	y��-H{Զ���v�	|���*Y�n,��`��ٶ�1�e��Zx�%�H�?�R�w���B���T�e������]��Bb	�y�.��B���)�[���1�����y<�����7C���9�61AДg>��?�w}Z��]�"l~�y���u]��Y�&/�n`=�L�<s���4�uz`����ے?�jC�P��֖�uW@5�UX��{���?qʛ�C���7h.(h�\
2q�̃-�i2LO���[�y �l�C�z��U�/�^^L��>%�1O,���m8|ս�)X6� ��{�Uf��cw��3H��(ֻ�w?���o���"8�o��Ǧ>��Jf!睹��gu�^�.�;%��2�}��߅|D2�4�ӑ,]��X�����PՋ���ym؛��Ǹ����M���זI��-�o�Do�������O&u�A��S^A�M�TAa�rp���@�oқcHi���Opq�64�S��8�0{C�T�������7�U�IA�c(��N��m����������O�a�ZK(a��z���Q��@�7����)E���)R<c	���5�h� �uK@[�G;]O���9H�`K��;b4���t�35�l��X���kA�w����!k�S�`|���N ��*���eƉ���#Q�!�(T�2x�=�o��#7�����Zr��y��k�D�$m5�Yj��G;ҹ�K�n�z�^X�6�ӛ몗ďZd�WD��R]�[�����f?[�+̋r>C��DN:P��Mo�*2�̀1A�:�N�*ETR��xſ�Cֲ~�+�u�-�%�C���o��ʉ�ڑL����Û>]w�T����m#׮S�3I�u4xx-xb1���X�@��ƒb3��#���O%����7�E�x4DY�Ϙ(qH�y+خYn�ױ��1��	���u1�3��.A<N�a<������gx(����Z���q�E���5{��k�6�AF�1�^(� rΫo*���y�W|��Z8f�Bf` њ�+�~,<r;�����nN���AZ�2,�1�a|��S~y7�F��@�R,Y�U�Aȥ�!?^K��)��m����xkGn���/�H�Bz�.���J�Fm��x���¼�hǥ�|�A%��U�Q��1̺"j�8��#)�� �;JTƬ�9�F�Ȼ}A�Ex��ݱ�SspJ����-��<2���~u�x]�(#?5W� �z�1��wF��v��1�����7��lf��[6IA1�����#�"��}���R9�=>g6i}3�����Z�ze?���Lt���Rjk��C�i''ZE�ަ���w(ۉk!����״c��y�/7t|���Oi̐e�;v�*��g0/�_*����t�;az����;�zY.�&O]7��Ӏ-���ZG�``n�������H[���\It�M�tYAO���wT*6r1������u7���%�V 8� No���=� yL1pP�	#cތ)�*��C�k?�e�J��6��Tz��?>���^�@��҂�Z�"�.ʟl����7�����@��>k$E�Y&�I[N��n��n}+,�e&���IY����(G�`�d:w($�_�g�Õ��V�׮�V�� ƒ⭫`�#�r,���EPOLE�+�E>�T��S�p��ڑCx���ȒN|��q�j��`������b]6��38%�~r����V�WQ�g�~$�m���ڿJ��K��$���� 2����}a�8��O$��Rܡ��MS���uD$�kW�v�Ԫr좈�"XSl�o��緒>5�wkէnG���T�2Rйضu�T!_��I��h.�kp��S[���j�H�e��'�ug�����ͷ�pΪ`8�����-\#P=Ćgp5M�@'�@^�5�5�3,E��3��&�Xboh��/G�n�al��!���
��a����P&K�9ns����$÷	nܞ���C*��⇤�ݪ�rP��T��� �䛸!�1ܬ���2d�v��J)���Xsv�R��,g��e� �e��S]]�9xlU�:D��͗�c�&W�S�[���F�:�̙TW")t�/� �z�%R�ϑ#�bл���>�'z�����S���^{�h���2����(�x��:�\J��\�!T�̇FƦ����	��'�?(g�Pz��a��}Q\��=�/I<cK+�����E�8��SxH��AcQ�ց�Wڵd��O���t�\R�h��L+<Kl���]Ť�?|�����gma<S9�W2�/�Qo5b%���w�,��7��^HA�e&�S'��VeԎv�`#D���*��8Jt�d�:4�I�}SMV�\;R(=PO���&>�B�w\��_�w2:~a!�d��1"�8�"	A�+9hW�b,�N8������K�"Wt<w�C��"�MBǽ6��l~r:F�(%��?[o:�o��p�t<z%���n���h[�z�bBr�����Uݖ䇥�(;�ߊ��� �Z�]�?�����"�0�#�ʪD=�F�+��.2�� ����RC*�mA��>�b��Y_ȕ3�b��RI��,J�Շ)E8	��M�Y+�l'�S����	3�zn�A��
�澪�w(�Va��Q$pm�͸ �Urt��*�%��z\�����QƝ."�ۛ����/1eտ�	�^C�`F�P\��B�@��Ԉ���D�+1%�U�cA&*�R��Ԅ�ySP��!��TW��ΈJw/x�*�Niffzp��xY���j��yp^x[d��U���Pfm�$~<	����TkA�����1�k�N�^饴�����@I��cxLW�z�;�:�V����&�-U�Sɋ$2�E����Pu����Q��v��ޫ�hk׏}�w��E��`�#���x��u�t�;
*6N^�=*���a�=���\��t+z��`l��I������0����.9������ډ�d*-��.�ϐ�!p��^��E���F��{#���j�@vS1���ҧ����H󶟌H����:��c]e�'Y��`���@ZQ0s!�n>�w�׵:�ݲ�&\r퓕����z��X�ɏ̚Q���yZ260J���dEU4������N<_��H\�LOv/�@�?���E��89�dm���$sڍ�6�ڍ�~����'ʞ����2���r+g/����BC����
IE���$iR.�m����DC6�I�
�Nz�K��n�����Ct���V7Ҹ����3H.u�5-����`����$�5d���qp��U�F��k�nwS8g!�=�U�a�ѡ]��������n�yY�Ѿ�6�ܴS��~kW�٠��B��>��W�/&����k]�D�5߅�`J�A~���:;ᴹSUEi�ۓ�Z��Sg��Y�Rw�wG�kM�qT����2�R�8ӄX�hߘh�y�_�m�~�'�xf~pݑk��G�o%vzlH����t�o\��r"%f���2��#O�ϴu���$�CD��+�D�݈m���Do�<���m��ܹo^�kDfpw���#G<�hf�Ik��ؖ�B�������nFϣA�lm���DYa�������~�m�8Ð?�8�Uw4�v�n=3[�t�����v"�e^t7�Ge�B�c�ܠ�x��:�O���Ǩ��y�M�v�?4��� Z@@[<���ք)���f�G�1t�s���R���yץ9
�꘦>+/J`�M�Ҭ2JK9}sJ���yPݘِ�Iݔl�=��S�!�9'���c1��"p�`!U����j�K�}�T��Ɲ���_/�k ����G��:Ȭ[7������ʗ}�S�e��<�_��o�.��,���h��8�k��,#������c�s0 Ґo�A���l��&�C�
0"�|s�H��+^	��ð��L�A+,))�閝iZ�ొ[+��1�T�Ym�ٴ��s�I6������ѕR
����[2ut�l(6�;��� t$�?$ezN���_��4���[��d6'��n/W�Ժ�wƛ$��=& ��f%%uSl�ھ�raQ35�K�l�g��v��r��"kt̲x�D˜�+89%�ke�<���2o^���j`��9��rg�i�_HҤ�p)�Ԡ���-�{.�k��;�첱���XU�W�9v��M�Md������DJ�Ѹ���UҦdM_U���B�u~�[]�ˈ�U�Y�>���A�`�2n|�2�����uIsTN����Ba'<����s�$|C�� �>�bP݈{������n�l��;N7s�o�"�s82�Mݑ�5sd`��B(FD��T�X!Q�uƄ�H׵Wɩ*���[\�{���6_�
ݰ�"/S0��~D!�7/kS!��- tHH�Ƨ�/1� v
I]������e�`d�m�~�����I���D�X"R��H_L�ء��n(�|���sY���e'/���|e�H[�û���O Ҷ،�+m1I��ʐ�j����4�-y}ǟ��$]��O����RR9{5�	�8���u�C�60��3�I;n�HG��v���O
������8iJ>,y�������"Jk1km�?�2��m��������[�>TZM�I�b��%�y��<�4�@�kͮ��֠�Ը���WW���}� ��nͨ ��s���E��a�v;O���t�B&�[���W!F�|02٥z]��N�� ���ejE��K^N�tm�"Ac���p4��l��JB�?o*��,q1�$nTI��]|�ʳ�P5iK0{Y8��wT.Az�e9������	e�UP�A���s:��tk|��+]�S�Y�5�yU�L�.�:�]Um 8b?����qs����I�����'6,�v�3��Dc���u �k/���S-ĂAз���_���y_�H8H�I���5�s�T� �{L������~�xe^߇���3۠G<)�B�+��m1^�U�W��N��ND�-	ႅ�e�L�X�ʞ�O.�/��:��s���{j*�IL�*Iw,Mt+�5)�,��	�~7��ڰ�s����f���7E���G���bfZ�nSg��.��_˅�x���X4h�Կ��U�;��na�l8�<��8�<X��Nn����-�5]��j�g�����g����E�e���f�h��#�պ��O"�X��C�:�wR����8L��t�o,�X��L9��U٣�#���!�z����"�m��,���}�c񓩽EDa��S���ԭD��b��+u7[��Q����s�����l���c��Vq0eD|�/�-J<B5��85f�HCb�M�=@i�X;3����R?z���|�-+ˤs����ћ�US�u�ު��B��+�Y��Yt6/"��q�n&�!z�2<�<�$�3��H��$�������69E	���B���˅g��f�[�p�B_���a_�K��u
��ob��;Jd�����;��LZb)�V4X5��>���^��r�q�e��$��
T1��^?
W��G��oZ�CA�8}�l�Un�pH,8R;
:�˽�'�O:��Jo�F@���;�d�t���4 %�U�c	��F�((6���ri� �DğC$�z;�#.�c�2����H!P:�ֵ��
d4�)Z������*���������C�M�� �Bw�ķ���0b�4"$ًV��~�a,�~�K!����w#	.9�a=.9�Ǻ)�s�;+��		�#\e@|7S4�{���;	H�u�م$$��m����d�Ь������t�E ���v���8��t%C+��j�g��E/rUU�3w
@�p�l J����ঌ�\)CB��'%��}�<��A�]�C�ش��!��U)��.��hi	-��a��c|��ַWA!�9����燼A��{yW��ā��0�m�f���-��N�J�l<��@�Ն��g��WD�ɍ���I-��0�nS)l�⽁[:!	!����BDy�8a�y+���ٸ�(�7�-�kR�Ů9߄�]�k�J�()��[��r1�{؍)�3B���s��&4�����AZqypi�C���@^��_gğڼJ%�x�b�/��5?-e�V�� ��[��H%Er��lP���x�?�����0�����V�[j�ES��@�w�*��c�>&�$�GY���3�J��?��U���#F��S���d���k�l�_�z�^�'.Ϲ�}a4�
���/������E���έ����g �L�s{(�SZ��}x���N�2&fE�8N��ï�ɽ��7)�s�Y�����_�*��1���2#s(�&�?/ޱuK�!�4�y����7 ,=��X�X!������[�/_q�>�Q��0���B�_���,[�s�{In�Wȯ���8 "%2���l�QL�9J����tz�p%�j��G�_�ٗ:n<'������ɢ��RO.�C�)4���X�ɘ�ǢV��I<U/h�m�u(^FK��Ӡ�t��y�5�*|��i�No'���6>3H��ȾP�d�3%��^�#�iu�ܥq.=�V°)=4�w�vEJ��yy{��Q�Ux�R����9�u1�49nw����m��؊��L��lS��9�q�L7�8u�z+����޺�6>���|N��(e��}����i��m72��3R(��T
c,�����%$Z	��U[��b*���;.z�9�פ���'5B̩4SO,G�#�-,�y��vݜ�\+�C���Ԕ�K��PJ���!�C  �-����Rʽ
\Y��#�#���@T�qo=���7U�/��?;�	X5�粼j��WU�s!����Pzơ:� `/Р��Rޥ��q���:Dm��������b�j
��JLgX���Q��8�c¾��<�J�ҳ��VN�'i{ʿY�П�)Z��7��U�OG�����W�X;�ġqd
�?��%P7j~�Vp�Md��G�����Xc��!��L�G@�6����z�M�W\��Ҷ�كH!�2|��
c8D2l|���M��"�wh�7���5t��bAk�R��������e�}�R���-��伸[b n�8G���ƴr��;�QbʴmcC��u���z�XmtC���S�W
�@3�R8�׷w]�FW��*}���%����N���ǫGܓNt�Q��~\���E
�}���[��QKIVe��9bpq�c�5��1�s����R܊��f��(��r�㧆�E"�@]��鶽�<P�dg�
��o�}w��p�Eqi��:G�'|#�rM�ѣ�m%%�9�H=>��+�
����i�*%Htʨ~dB��)���XU"4�D(�fVϩ?�,�m�nu������	��_^��θ�¦Ʒ����Ӽ�ā����0�S�f��mJ�Wl���1��i��L>xn����L�T�X�l�G��O�.�N�3�䂶Z�KFQ���т5C翾�h��cM,b��0?���7]e�� ��k�;L����X^ʈ��>7\�b��Dpu�a�D%�4�����,�6j������eR�FI�`��Ǟ��J!H�h-������EU�E�MQh�ϻZ	4�b�/_�xtA�^����U'���+֘m �����2���K�$D����� HeC���sVeI�����2b��H�RM�Z���z�Q���haؽ� {cS�r��c����I[��JaUF��:���L�Y��t�I�$�����r�^����MB	S�8�A��$ Q���^C��P�7	�nf��F:�}n6Y$WP��y�Ȼˉ�订4Q{|љ���)皪��C�KX�7",Tu�s�V.䪾��E�z��-���d�՜�cީyW��hj'ƘO�o�� �Ƣ�+T	:� ��+�T^\ء�,X'��-��c7r�U��E�DR4��j�j��Fh���g�Q������{\z�ZU{I�U�u���S.�L�����l�ryʍ�oy�!����������Wy��X�����U@�K7��¼&�������_��o2w�Qz�Y[�,]W|W�9�5f��ts@�>��R�J�>h�?��O�bR�����þ�=����/�?�r�{L�_���WOC�����SR�yf��?��_�������ˇdw����K�#��5��=v��]8 ����yF�5���o��R��l�n�V7�'A���D��~������J�(��JQb��c�C��HP�.��aR��W�j���Lg�m+�ư�:���t$#���$�F�jY�����k
�ż@��ʚ�#'fM��1�o��������<��2� ��uE�#�����N����in��42J��e����v�v�x����|���2����
_���eE��ɨ�噄F`���r�.�HW����(>�=K �F�%���G�w�3���o8?�T7�����<�։3Ϝ��lh3�z�y��s�:�/�r]@Y�)N÷lA#;������Bd�f,����W=�`}�bi���@k������zQę�N�ژ�m:%(�,\$��`[UFP��C��
�> �h8�5?����V�d�ؔ�NTNAP��$��Q��Ԕ�kw��¤���������槱}�~=%!-��>I��_�RU"Y��a���6;���ВoO��)W�o��`{�1Z.�䩂��ٙY<�:����7;�f������0�0ֺW��I�L��3����.�=��DM�L�h�Ѹ�ϮaĬ�á�"�}'���S-�]��xs��b��տ=�Ɣ�l=
E�$�(:�S�k��MZߔz-s�.���u%a$��yE1��|-���Ӕ���>�h1]���Ir�Dl�e�7\{ �lyI�\gt-�ZX��Px��^��<���V#6Týtp���o�Jv2�~��5]*���\�'&�|���>ix{�(�o��R#��	���[��$i��a�ŵpZ��Kض:��wٕ�����	��T�v#�����i�%G��~����K�n��Έ��	�y�>���)��O��.>�N���IS�����?�S z״>��5Ta�ߑ��˘Fx��^Nʛh�$�HH�����-_���t��kzI8&�+s��om
��hX�Ǒ:kN���+ϞF�"|��->4��6��	\Y�:O�t�]��;�h�亵o���y2B$eឳ�~:�~8*�@�F8��l!�4�gS����?���ށ�J��~�+E�Z�������O�X�����L^S0���i&�K�"�X���
�KX�#��-�ɺ�;v}R�;	=��NUʏ\8z>^
�)��F�Q`�f}ZB��\'�]F�u����(� G���Ӏ'3=�'W
�` `'�0B�+��-?�#�S�ѵbf�̞�ؖ���Q�}��a�a#�*��|����"f�QZ����ęŌD��7�a�+j �ж�sb�X4͐��(�>��Af������q^�q�q=ai��!�x���Œ,�.��z_�}(�/�(�z��A��i:����.��Lh@Mf
�5�nΔ]Z�A��ܯ��E������H�+�i���S�H�ɚsh���x��d��&M,��8$�A0F�<���xKX��>��b3_�s�hz�ʦq���rW�%���Ȭ�t5���	�����u�~��qŲ�ˌm�mM���(�dP��un�S�pҍ",*=��b�
�(��S�m3 �Ҝ����1��34��q$9a��)'z*%S��rE�K*��E�W$���"M��ȍIڋ#_��og��sA�G�� �n�<�;���$�v\��Q�t�WM���)��XV����b�y����0l�)�mFz��s�9��L�%pI �	���O��-��|ۇ��~˴��ZƇ�O�>ڍ�D�޼^&�>��Wf��.6��yYP`���	��1/�N���	���������߮�������z3�[Z"���pg _Z/
P�BVQ�<$��R ��D��/5�PT'�T��<Ֆ�n=�\!�8XcFO���K�d*�f��,cP���K�WC�2��J�x�o7���r���T��~���?�Ϻy�l���2�2�5����U�	�$�����9����dJ�~�<�[ X^�#����Ư������i�����K����2�d�3�G��Ƒ˧�0��
2���SA�G�\Map� 4�H�<��(�[*��Q���̧,���D���� ��������ʷ���d�ʤtU�<G�Ƅ�����T�07�6���pH� 
u��۔�iX�&'�Ch��A(W�W��r��L&��탕V�L��/���-u[��ooȧ9.gɰH1��<Ӿ׀P�Iٝ2�'$���
�e؄d��R�����x܊��]~���j'3��U�V�s�_�.�<�=�����aQUyw�< Α��D�CNe=����$�����o�h�^xPc���:���Q��-\$�B-Ǣ����
5m��qc� ���a�%��ct�Ȩ�����{�-����n��o��M�Q/!�]g�h<3��Q��|.!���vw �g��=��Ek�j�(n��C�j��vEK���nڀ���KtЄM�b�iV�,ߧU&������G����b�E`I �8��S&������-�zS��(�D�+u�	�|��Ko*���#=-��a-��1?O�V�K��á�g�a��}C��3ܠ?Q+H��ߵ���S�~��Y�9�Ʀ�c����'���I/Hw#���� 'n��p#��<p��V��i������?/3�x =Zu��1(��Jex����^�`��_�R��N�QF�O�%�m�
�/!R�'�����;>P[����ݏp~O"�T���[$o�<=�9�ӆ^�l��[�zDNb﷌V9�
w��9{�#^m���\�#n��7�}D�m��f�&H�i�����.�!K$|[r͌b9�Yf/�b2�Lw��|]s³,<@�D>{�.k�,s����uhp}� &� ���e��d͞�^����G�\�Rb�\H�K�Ke���㺾����A�}>	פ�?��G��-|��o@���飒H�ݮ}�8
0`c��%�c ���8y��{
��&������x� �2��ɲ��6[��C����\�/�`�f�����"P+@�{dD���{r1޷��ߨ�s�`Kd� l������a����Z�г���R�eo",��� �t����~���M/�%,㶕�}+R���\�Sָc_�ٻ_�m8d���_1�d�C��V��v����M��d���e���˧B僯W�ǯ��,ZI��7 28�'�~��N�x�W������.oo�^�G?oRwʧ»G5=�c�o
�=QĖ(m�����v-��k���� �˰"cQ?|��W�PD���.���f!m�������+���&>�jd���T��F����]�Z�����t��R�)�)��3ݵN�qaȱ�릗�H,�� ��+
�2����FZ�v@���t6!W2������ P�n3���̸]�ǳ/�L��*�[�U5��e(��Ip�N�ve,��=��h�����|�^U@���J}��^5ƅ�+�'\H����[�DL�EA�wLU)h�0�{�X��M�e�6���ڃb�qk�-ޟ(:��
|��ꎡ���u����b^�d!H�Y1�ژ�Rj`Vnj�*b"*>B`cYD�2;~��|�h!���u�q���
Q���7��H�_A���lʳ�b�s�}J���n{W�q9��@%v�E�6�$��C�wG���~
Teltة�>�R��`a�?�~���I��ƪ�T�K�^1������������O����SU|�dZ-/������.Q��@/�GP>�&�L���QlU���D]�\,�	�������4��4A�J#ĭt�Wf����) ��G�<���"@ �:d���=�K[R�-��.�6N�`�Mx�䋿x̱�1�x�Ęr��n��~�.��~^�\A����`��AU���?N�Aٙw�S��f5ZP�Y;��#$��]tL�	4j��բT�6st�7��4�G�� *�m�Wsl�π�6�8al0�#����D`�{A��P�@.x7�S�����ݴ�~s�v{���h�\�lR�� ��,�'2�z��=�*��R�����F��y�^��˃+�F!�hE�ab�(y� ��kN)U�$�K,/c�OG��I],�hHbѻ�M��"�$�P	�O�:��Q&��;P�O�yW��0ژ��ʝG����di�����L�Io�^l���� }ie^�	<��?�m�	�[�4�X����ﴮm��+ޯ*3����ـ��:D|>��L-�z�h4r?�'nB̗�kؚ�v�bW��6b���H��0�uz����%�'Ҙhҥ	����c�"8p���
�r��k��Q*;�8'y:beĽ�5�m1f�297����2����� ���nZ�U�I{��0**��ar�7�Ҙ\( ���Ԑ#RS���c�f������������Y Ԟ�Tz5���C�S5N	�>�-]X<c����PJ���Mx]&��B�vy]��-q�Г"?�X���[���e�IP�;�<PNm�yh]�*�9 N��_h>���Oɣ��Ƅ/���Epu�o:M����O��8�.7�r��?	m'�t���c{m�-�cN|Ӏڧ��u��G�c��ҫ�E��+���!e�ˏ�v\�r���9*�R���7"�-f��G��ꪾ��W�j��c���n�^�&8O����v̢�9%ם����m6��
��,�4���l/�^�Dx�ٛ���*'W���	�E3��C�_x��}�Uvt{����%���mN�\	�ˉKw�B43	?�/Lku%f�a?�e��b��иl_5t��/fw{a���`�|���৭�@���H>��
�3
E��;j�o���)o��'�Q�+,�r���@B�G5�s�`)~/a�s&����Ʌt���45t�8��"wF+ZS�3����C^����B�&�X�o4�|�jo�Jqݕb�$ׯՂm��e<@dOPK��8C�'������	�jܹ')Q���й���U�U����t6�S$�r)i�!��q�0�=Ɠ��A�Xױ^!?��73�s���(���� 0��M�6ͭ����f�������.����P]]_�y���j�roj#Aؕ�#���ش�n߉��-��Q6�� ~PL5m��ˑ[.&o��L3!��+j\��!�VL�㋨Yu�ؐnl 9f
h�`�nL�����?�qWnkZp�&�'ʹL���@�1���F��L@���a.�Jz~�a;������8&���, X�����p��z��FQH�7V�ֹ�p��Cːl�L��sS���/pC�Cw�}�2�]pn`�q#B'l�֕s�H�M{�(�^�_�2�u�^���@YQI����alf-����!���EF��T��������ml�ˈX��}��plk�lmc�*.x��{��+(a�R%�<�H3a&=�?�hr���Q����_d]�sp ��g��vK=|2��+��y�\$<-Y��C�cԌ���]׵V!�d���4t"��l�$P]v��Ã�S|�;��u��	1Ws��Jݖ!�B�36+�!�D�ﶜpiS�Q��f�dqV���q����A�L��k��Z��4(;m�]0�,�����/�fP�µe� i�K�)��\�D�3�8Z����'c���,�#�}��>ΑɭH�:��v�4$�Ɨ��6l���c.1ߪ��F>�w��"	����񘙭�r��{1�a��qa&�vX�"�v��S5�����o�̻��|T	�h~�����3q@4�0i4lKݓt����앙�;-t�})`E2��+��D-T\!b<�@:L�I��Y��nl�G��-�A&��,�r6��>B��`��J��bކ��>�kQ��K5�{�]�� ��}Mწ���ҺɚzC�l�߫�4���M�yϠU��n?V��H4��r��xfml'	K٤��){p!	���{��Һ{����Bt�����v��.��n��2-ĸ�^	�Lw�{f��Za�gFX,;��ugjnm�մ�+4lػ�B�� O%tY����:L��5i@SHR`c�9�� L�,5䈣;j��nk��'�i&����E��4�rBV�'�����d�� �Q���<��I\�2{ߩ�9 1���]�Q0�b�	�����ݜq��<�Ӥ5F�)����j�j9/*��ߎ]:�^<�:�^�W��O���U���(g�/�505j��c�,X9���χ�Bb�I���f�hct�	˞Z��{�R)�Xz&jM�E����5���B�3�j��&x^��ݝ�l"fZ��I��U�,�v�^�]���pL<�$m�v'͖�C<Aχ\�yd�M�%�$�G�͢�C�5��k��[�B�6���֗�l�/�3Cfi��˕�X}�H��	^�:����ḙ��ܪ��1g%w�ԁ_���|+.�;E]L���nk	r�d�'�F ��(��<U6c��Pӎ�d�Ϝ~f���h(/���X���A�W�����]sءJ�G�3@�J}��s�ŵ�h�2�1��s��ʌ�jyfK���+�|�D�A���v-�E�u]������YGE@
zl�g>Q�H�<�/����(yY^V�vV"�~�T��A'�c�� ��r�O�r��1X׾�6�FVu7�"`*E�B؉��9Cp�-_�h6	J�_��M\�g�$rA�1Nx��M�QA0�T���bj-y��ǅR�@TI�ə����O��X9;U��3�&
lu�F�F}L�Vuδ��x:�r\;���XVD�>ߘ���=�J ����w�����u2_�гў��#�
B��;�[�:4:U�� �b@��<8�����&za�gFI��:�
�V�%K����1���5�9'�
�G���ͬ�"h#��|�H�ݳ��'��d5qR��?YQ}ss��N�����7��PG|o��7��_��p��۽|���� (q����&�6%�5*�P�@R�\�;����d�raY.�iy��㻞6��
HD:mϦw���(����o&������̮:a�G�����b�ߤ�,�J���P�q��E>�Ϫ*DxRQ.��B���o
�|�]U�נi��9��*V1��zf[�v�
F��Vy�ؖ�qnR�б\Z��\jb�U���:���^�S-�D�
���d7��hH�;�k���UHշ�%�|�O1�\IM{��T`G����<�'�/��o]����Pv���Φԋ9p�����?�K']���]�i�X�e��̀��>�_߂���7;�ܞ�ٞf?��Ja��|�@s���3�=�)?����,�lI���ޗ�Y/M#�13�$��˧9���m���1�=�v���m�`L�JD�1��>Z<��)�?�m�2AT?���2O�?�Iې�2uQ�$:f��]ţ�$������.8R���|�S�����̹���W���~p��8�	�Pxj0�j�糿ה�12��KT2q�	��5�Gp��1)�ן��3kEך�"*"l�R�U>�a��8��!�Z6��+��[0��ٛBQLƯ_8�Ot�IH5+�<jY���M�w������I��L�:�c�iHa��3j?(�#q3� *;��d%Fd�Xm'�	�'Ƚq@0]�]�~��"��y#��2WI��UE?f����"�x�4����K��4�$ʐ�O?��Ӯ�c��-����԰G���3<��XLOl�-bQ:�p��.����s����7a�?v>Dn	����ew���l���1�Z���*|����7t&�sr�yy~Շ�&tE�1SL��FxxD�yN����#���7@*�tgLCO���[��@w�^�[S^h����y>^)�V�|�@~��{����s�s�&�E}�W�h�r-78~��8�?H�s���s��÷+L�c~��	r�Д��xNH;=�wO��.�)��ч�� ���J�ɂ��^0�zM_d�[��&����>�K�j�`j�!aՇ��FT#�hvQ�ׂÄ��o�ǚ��.Rmо(��@�(�L���K6[�(տ��%T�R1�G_�#��>4lD LT��2�$?E�N�s�|�#$�
G`�{kcA7�G�w(�#�45����Շu'��έ�B!	���71�xz86�y��J'_����>�e�3`E�$�|�<�WV]A�V��O����]-�*;2�:�����]X���OI���|�����y
�@���s��jN�j��1��� ��e�:�פ0c�7s�O�-5O_kN�*�rT^N'����U�ɮ�V��u�]11�������v-h~*
p������<�����ֈs3Ex����S)5�*S�R#C�N�1���%�V�y�kQ ���}�TE�D����8�����53HӦE��5}��?��E�>h����q,�c�Q��K��cE�y�:�'I�W�l���Ӱ	==)��ԍ;e��u��E�OE�e������`���zIR�b 齝�_ϐ��T�Q�f����um�+�*�{!�� �M����.3:Z�u��,�Z��'�>k9ZS7m��ׁ��,7S�j�[(�Y��6D(�2�\&��KM U�u����1$R�{`L<��F�����z��a�|�qa"��،��Y�f���iZe�����=��`���7,�N�Q,���/�r���ݎF�.U�=���&��y����߻�]n�}.�3�v4<4�0�5��_��*-R#�V��c��w�j�v�����$�٪�ȟ$����߄�0�#���`�{�E��f��1WhI|�˗��1��F���8cs;ʭ]�GU�O`�v�(,c8n$T�R֪�T�
��Z���b��_�Mק{㽝>-��F�#�,8�U�ݜ5F��]7GS�4�������3|O]j9�4HS��1�)CA�e(�h�E����ޙj@r=���$��`B�RPݱ�Ѐ����4�x=�O0�Å��r���Īoo;�O�R�/��x1~l�ϡ#��ʜ����}ok���/�t�~6=�n�5��Y�h��w�� ��F٩>�j�:��?*D��,o�}�#uMDɮ@hvH��&��};�9���l/ޙ6}�K<��^�V��.�Z�j�kA��X�/�Ǜ�����Ɨ.)���/��� �${�H�iϬ�<X�r/�}\��Y� :m��qAN�8'R`� �̖�b
�z_G������ «B�X�	7���L��/M��#'��3mҜNq��mod;WP��w�o;n�̠�7(��k�묣��үY6�Za�_� �Ą;YL��w7!g$.�:.�+�2���|����t�4q�6Y5�qq����A��9�l�T��m�@��cl=�e,8��q|�o�|��o����i7���P�C^���|`xK��'/�A��6�#^�q[��?.xx6�)tgT���щ�\�u^���[W�t�\`����9Dʴ�4��!��%����5�"`�x�����X�YhE�9��K��[�#DFnU|�=��U�FnpT�3J~ q��<�w +oy@	k���ͻ<k�����������	� �T��-ȟC��"�ɻ\=qŅ[~~i��y����O.$;���%&�'��]���e��)���%6���
�߾3�*�p���w��&�+I���㨲��jzq�fkS�<~���z/�ww����G��_R�8%P��	�5����F ����5(]��_�l)�p��3����(�t�B�my�X�Ts���L������	�b�Y��;8��Ή���<E�<�C\&cOZY�U��+�i��vL�Ԕ���2%s��O�+*v���H�8_�Q���%ߛ.���G�i��T�z���>������;�ypd�t@=�h�J�Z�*�B��p)|�̍_�!�����p�.s+ R��%%���32����ei�<��3ꨢT�_ʋ�\������^��Bn��)�r�L����/�:,!�Uͼ���?�i�X(��Z��C��N��Q؝�
b_o���^@�G��b%
%������ ��f�1���t5�J�S�l�;���u�$~��v��>�c �����rw3��Y�:*˸a��ڇ�;ȯ�8'8]�Gj�ܨK��ӭ���0!�H1��0^ky���-G�2l�מ6�t��e��Q��-��y*�̮�D�B�CԚE���Pڞ���;n�O�Zi�ϡ4�C�����sI�& ڴ:J���}��l�i�'�L�Ww>������5�u��)�?��]�OC#z6�;NM��u���ʱ� ��ky��s�qN�;)Lv��O������qC���jsMFʸF6������nN'�ܞ��?w�j�(���0�p�*J M�?�����S��j�y�[>:�Ű;lh�?8Dءms�̫Z��MX���"������f1���㈡|�v!��e�iR�!��z��9�Z*׿kP�f�@�lyK�v��-+Um�h+��s�� �H���T���d�TK�zS	�`���ӻ�'^�ү҅4�L> K����zYpt��sÍ؎�
�Y��8��Y���X%b&�<Bط����x�Q&�h��LڀPh�I��S0PY���S�=���W {�t&���X�")s�BU�t;kcN�ei�ۡ��aƤ��c ��.��H����e�H���(�<d�[��g� ;j�S��<�pպ=����6�$����u�Is�'K�vuY���
�Ծ
N�9�IOqK<��dO�6D�%���*�;�����̧����Ő���5V��
ZV��bL�lQh�ٻ�#%/�R��a�t�����8�~����FZM�;���H��> X�d"�Z<���	kvj C�4^ 7���w�����6�e�S�4-��Gp����Tr$[��~�&�K�<�����m6^sܝ�.�m!����acQXl��ƛBWW& ��q�q�  ���i��_���sg��c�'L�1l���'����L��6OT�ʜ�����V>O�\�dq��d�iv�%n6$���	�%]3}�TQPk��ģ�^� :���F���^[�.�� fΓwI���H����e��7���x"��HA���2���O��Y+Xw��\S�>����i0yrr�A:긪�)vp~���M8S�|�wXIJ�Kܫ�{܎�ʜ�Q�i*ք`�{��J�O�J�,�D"{83
;ۂ�V�S�x�}p|�zx)z��շM����GE��ο�]Q�P����WYpt2�A��
��Ad��ۈLZ���3^�V���op:�'��N
��|�9#s����egv ��@�<Z���n�*�L0��b�I���~0��U����4e.��b�O���9�X����ï�?�V'-Uu�K|���@%�^(_�&�`"m���Ca��W�;�zmm����1���*-�뢩�+��i4�4e�k�r���A�e^�����9b+#K+��ދ�v����MnL~�ǇHTx��܎"�~&pe�}˧�Q�%�@5��h��DK6�B��J��<�ݿ+�?��,���[��?���lF3��K�}���+zT�qfv�J,�\���{3�Ha�)�/A�t�$;X��?�'�F�"���7k?�D;ƾ��>x�S`�#���pB�+Bģu?v,�)������QE�?��Aa��g��u	c�/��ye�>�Hun�|��"���=gſ�z=�Ɠ��=��Zi��A�=g��A�J��2}<�@��B���F�oPK�P�L�D�p���)t�Y�9 G[S����K`v�����T8��)��Q̊��[0��^�#�A<dg�ȵ+�!��7A�	G8b5����ʘ�҂��u�	�e��A��&e��c��Ŷ�l����zp��|k�J>,����K:z,���۳�R��O'a��7-�	�f���Po�n��[����Z-iR��G{��˄ 5*}��s��%���*���"Ff�d�Q�O���@�su����1,�N���A#�S���+}��8�b�>U���X _6���QaT�g�5fD���H8�������y�8�VP��D�kX�,��Ņ�Ć�!N\8k�w+X�5�C�����.���j�ŵC(D�U��$v4���I�ܧ�A�����C�6���6�Z޼�YD��]B����v�t�A���宻�L�M$����9Əy��ȈEF�݊ @�}7�.SS�ț�$��0τ�'=c�y��G�hViy�1�7�:g��%o��}�1��Pe�ox�:���^��7"%¦���� �RK��Զ���;i���� -��Gd�H�uW(�?+{`�ffr<,w=��>E����K��I⬃��AA�++�l��{�Sۃ7]N�<K��?��[��ޓ���`���,�����ʰ�q�ln�Q�%�xr��瑼aʿ�aN��=r#Xٮ-������3�zd�L�6=iA��S����CӔ+�#��_v�&+	�<	f��C|�0���`blmO�6R�r���fS�]�o&5ot��Aq��,|� m��=e��%��z�ۜި���v�����x����'��&��Z4V��;��z��y&KTi��86{����RMCW�e ��pkPzvN�lP�6!Z],[�y-��O�ZsK���7����krMa���� �<�+ލ�0�{ه����\�R6yz�t��j���,�*�-��	PCP����޷&������t�'֦։78��G���K�}�M��c.H�(�'g$�S��d��֑���^�_̻���[�M[�9�hݬ�?a߄�c�wLNG\.c�]$x~�oY؎5LR�H��83	���&��ɶ������[�rd�����W�/[Cy��<����~�/�91~�J��$Y0zVd�%�2��2UАsi�8F݂G��ߐ��a�e�G����ےmZһ/V���4�(�߫�Xe-G	8t�3ۓX1�&f�n���k� os*2�/��r�v� �Q�RS��/�w���\��%Q�;3`�Uy���3�*Y���Ə�{bRC�=��
e4$CeȊ]Q�@����C��\� i�wa�-��?����ͳ�:��TѰ�� �Ċ7�G��X�2+��%:��V�4gJ��<��mϮ�Q
M��l�����i�v��h��8=kU�b�]��DڽԖrd�3���Wª*�pV�eU@px���n� S6h\��gC8��Y���z%��4},pE�p�G�<������Cs.�Pfea8��K�A�
���*���-���fXA/��Z,��x�|�E�3n37KO��T�8Uޱ���	lA죪�#ʅ4��n��ñ�7��eh��Xo�ym�3�����S�tb���mS���M�Y�����L~y�^�v��zp��3q��RP&�y��-��:��������x�o�b���jlE6!2T�w�����pJwd��Dba�F.Rwf���Be����q��z�n������K���7h�,{�������	�#n	��]��O�P#����_�ҜVO0�����5Xu�e`�\n���Y8���?��`�����U�b��w�3!7�I-��4�����N���;�3��E��c6:,���.�a���.��R�O��_q�W4�����/f���Z�0��ɻ�a1�����ϕz׫??mK�$壕��p{�	;�b))�AǷ���PS�������~0� ������c_νF�{�3lt�M>�q��Qr�Ӗ�A���j��
d��1�2�#S_�C����E���%��%P����:�i��c�9y C�!�n����&イJa~�s�� �e�~|��0�DY(n�����'��x�Lj||�H�.�r� ��^o�Ƈ��:��e&a�~xVT~�"X�ދ�K�|b8�+{&=_Uβ�+I�%Ժhm�ҽ��Fh�^�A��
�vA�)� ��fN+)�������U=Q�Nu���#���h��7���}���"덥Ч�0{z��0�jA !�?�3,/0�Ȧ}ӥO��V�,t�ԟԤ;u%s�c/�*� L����������d"܇�F3X�T,����s[j��V�aS�`��:�����k�Ǆ��;�Lh�J08q�7�R�
����4h?ŀN�NzJ��^A$x��^I�M��Q�T�w�O+�j3A4���S�m	8��H#�P�<.�_�R�֝��vr��	�x�h4�P�%��kPVA�b�#�moڱa}��Pv>��+;ִGLK�j5�����*n][���Ȏ<��[��<�����q'�#����Y�E��)�5��
��(����>��N��	x�cT�͔�t���6q��m��L��7r�2'��+�?p^Az2H�0�ؐN�!����E������"[09�v���蚊�H�� �E[�VR�������$�a��*M�L�����Iժv�����@�R�*|uT7�؛�ؠ�Z�٥������I�kѱWZ]����)pm���|8ε�V&�S컴�,����\�{�:����oW9@�������� �
���C#X�C�N�;��	p7��A[���f�U<�c���go�p���>�����W}�&j��nà{��kV^�Og�4\Td{ JA��{�OF>��x�����g�cɅ0m3�%L���fU���w��8��,>�r��o���ڣ[�Dړ��И5F96��3zگ��x��2#����TQ���	R�_�D�w����*��� @�Do��Ǡ��J�hW�n�K^ �}4Ŭ�
��fd6�K�l#v�U�*ɺ ��w���l�.����d��h�<f����3�e�01ӥ���P����!�8>K�-U�ԧH��TH��?�N頳��ɥ{ ����ÃD�5��8f-ZS�@D� a�
�Ef�r~�w%S���NМ��t+��V�1�W�J�x����A?�Xe˵߮jr�uz��Z�� :ZX�q	^�ᚓ��\>�t���[C��Uo��Ð,u�}bV.�A��`'��L�^'���5	���b
#�,˫�:,�Љ*�/c*��yw��[m�T)F�ky1��HART�lD�x���Hn���*`���^��=!�.�#�p�ݙTS��(��Y���5�o�/d��Vr�wХ�j� ��jo�R��"���	���Rg3ժ�y�����Q��R�(^��	~�a�5��8r���%,��`�(,gz�R�-�!�a�d7+��FS��(�tڛ��[X���gA��̂��̶n��ȥ�O���sGFI1C���s1������e���kp��Ɏ��{j[�0������!�e=�(z^H��eR�B����qzec>>h��e��O��U+*-�!�{lVa������Bb������j��Ȱ�ϝ8����6��⥜r&a ��e�`�b�ݦ{��A����� )u���o1��ڊ���ri��ԟaZ�FJ�t�p��q�AU��&�@N/Z淙�ɻ�[�?y�Z��������${y9��}l���ó#dQ[�..��<ݿ���(�ص"�złS�Trr��5�����,�wļ��HƂ��w�$m� �ǥW����U��U�H&:�?@;v)b�bu�>N|?��О�.ln�%(q�G!K෣k"nC4�EDb���x����A�n}7�Ug�s��-`qYL�n�=Dٟ� HN	:��"�1�6��`=\�}v.f���P����`�1tղ?c��e�(M#w�/�
n4
J�w��Up��qD���&Sԇb����!�D ^��m<�q�]�q9���U�����%��7��{��/%�:�,�O5��G2z�Wb��<Q�������#e{�T�º����s�i���A�4�N�r�+?��B�J$�:_��^ѣ����s��2e��EMo�*A��|�7G�@[�Zoc�Ű��y��T�g�(�-�/E~� i ��rݮ��Ӹ9$�C�,�Ϗ	�YC2N�7��`3�V��1��L�8�,E�#$�b"�ePf��3j����P��\@���FK�g��`_.�e�*��^|]:����)O�bTQ�ĜF��[�l�u���,wxe�T����aZxB�-����[�A��V��=��w׊/Ӯ�\�������Zx%�Ð!'�i�G����Sy~L�Bݎ��ً;����ȥ�*cs�/i�H�)9q�1���l�[`�&�g�9�뇚��g����6�S�:��������?�b~���	����c�g��W�����^w�SQdQq���v�UwT��n��0�����x��?u�H��v�;���3��S�ʠ�w=��օ��Q���[����) �*��N��F^��f=��@�Ey��.��ok��<S�|���\�q��y�����Mѷ�1O���zM
�%�j�U�>/}zoG!+����u9(
j6�Z扨n����2�+�G��@z����40��~*U���sK�+�K �EW��P�xӲ�M�?�6�<UU���V]rbG������(
YqZ��U|��J���*e��mC����ij�i���O@��d>K���>�-��o�%ao�ny��c�D����wI��۪�ʽ(�#E��d֖��*���Y�
i0��Bi�}��Ai�Y-c�G!�K�:̟�R1��f��6����y˗�,���pf�ʢk�?Ԩ��Gi�i�U!t{��t&�q?8`Y�t�T} _�vh5ҿX�,A����wn:���tz��ջkHL�H�Ǫq�<Ё
P}�y'kу��L��q'E�;�OB%��ʋ�ѐ���-�1\ւ��7J>��+D:��(�Y)��U!J)�kЍ1Ǟ�/��v�f���a��5���g�𲙻�[�%�RJ"}��T�AY�XM�B�G�	),�pm���X�EX���5�^�T��G����^��Y��7��g��1�r,N�i1�~(��|%��\�6����c�}�����?�����q4��	�V���t��Vf����yW�rՅ��X��˪��wG$����Ϲ��?u}�w9�o֭�>?	bH ���m:0��Ud]�[sƌ��?�_�0���a>����Hy ����[.����Ia�i�Bq���e"���sP�����"8Y�i�\&J/\���+�5�
��y��mW���Z�?� 2��93LI�ڣ�l|g��t�S";e󚎱I�fG��w7!���6M�0Z���Ny�^_c��A"�VNq!���)��ѣn�f\VB����mF>@}F��e�;`��N�QO�~����ǲ���/����_��!%�_x��0J�F#%ɂ���J6N�ۇa'��Y�&<��qB�p�%ΣOq���K�/n-\8���x�l�=�s�s-��w��rДޅ���}E�L��'S�Ֆ4ӭ�؛H
�ںy���1XFB��=s(NTP�0Y75:O=ԪbRI���bj�m�n���IU�Bv�OY��\P�@��rʥ�jy��9� ��<��W7}R6�U�=���,�x�!9r��i`y��%��T�7��@N�����Cy��S P�
���TV��z�V�B��I�٪�%��(' .��&("W���{h�r22>���� �̟G����Fw�+�����0��
DS�"S�:��H2vï�E nmh��J�jG������%=YЋ��)��G�+���7��P��� ���	��y�AJ�h���bp���6ŉV�� �r��ٺ%�Q�˥�gT���2,1���|M"yO��hvu�uo~��4�6��R����i	��Ƭ@*4jmH��&��g�,:���NJ��O���z`�nV����+_��/ K�p��ָ��V6����qz�+$%ZK���T=#�
��L(r�`��E���Z7$�|�1��.�%��@�):����ԜZ�䏲�[�����g���Md��9��gip8,g��C�h�A�?�y��̫�a�ot���(��ݺ�F#�ї��<��({	�E���!��e�u�B|M�V��[�C-�yL�e�Վ������A5�ii��ʛ�C]���G��]2�4*}ԦdAu1=��l�`T���2�Ǚ����+� /iXkG��h���+ش&�6	-��/00(�Đւ�3�ÍZ����8��ץM�%:��FJV���ȷ�_��;̭�#-����Q|�^^�@q�࿦��`�{��I��T��C�##��Գ�D��$���H��CA寶��5�`s�8���F��a�B'��|ĢrJ�����h+�PK�-���Q�*B2�fd��[m�}�L�i����(�%�wT���<C��>�.d̓����ihI�,w��T��٬\S�$n�_}�cyG�)&��9K�9���b��ӗMԖ��>�o`��)�D�����@��"ŏ��$ `�For�]�+�D8=?¢� w@R�)U<�~Ǩ�.X�щ �x�y�?�������fǋWw�,I#��9�:]4>�QI�u��tj��ئ�ע�l�T��z�w��H�<;f�W�c8 reM΢�@�9��������#����:�Q�kO
����{]��P��:����YP�ð���q&K�Bw����mD���2�I�f�yʵ|�����]�Z�^���!J�d�_��lQ�V�JE������P ��É����e�	�(T���x_��U��i�B�\�:��V�`<�����^�����{ZG��6�=o�-'���-h�ٹ�����o�A�+�z�]$�"%�;s;��8n� ��o�D�K]1��y0u
�]]�̲Q��_i�������v����dq�d��l.�{��%�cjr���v��zw�����!�G�ýX�$�%�c����S̝:�O�.Q�k�PZ�@�#�~Tؑ�B���A!��@��K�~�I5��t�W���-��_��	χY4+�LVo~��9q�ƪu�pv�Yy�!��/�ը��x:L&R/���J�{9pyU���<B����+���ꍠ��z���>aUh@���Ԥ�@4 ��$ݪ���3�������5���=�K9l����l6�ʛ���њx��F�,�s���M@>
=�v�tM��^���̩�E��j53iŅ8�|:ٝ"Xi��&�FMI�(���}������,����n��˴d�mv��:������_W�!�fN�Q(
w"@ٴ .�IԞKf4�`�+O^�Y�0�Ŋ=��}�nG�b"���<��%��uerT�aC8�l0@���	4�/FR1�j�s�M	 %o㨄M�@�6�P�gږ��@>�v�FIDXl����&!�A4Hq�f{����a��﫭Ԙ��$ʙ�ջsV�Fd���k�T�5�r�?�H_=	y?Z�-_bnׁa�7\O�^��l"�m{�3f�y��2��7��=XVЦ\��������3�t<�<�w4ʳ+D�+��̢0�B!5���F	���H�B�yٰ��c�Tg�}Uճp>��������L$�4 ,xcH���r  ��$ ;/�f�K��X�6����t��#^��p�Yo�)?A�q�$X�A���<���V��DLԔ�.m�>��a]�ê�!z��0!��/��f�+ʀ���7�F�X�:8Ț.��8��9K�<��e��z`��p,R��<߿�>+�x�k���QL�^�����R06#u���
�vF��5�{h(�y�%�2t�7f�[=�s���ol�r�!��x�O����:�)����LJ۽�mnME���5Db�թ����ސo����k�%dF�LW�����1�\c<L4}f��IZ��(u��Z��yN����K���4�����6�(�83Tz����B��I�)3U���xv��`���?�����hn	��9�(�Ԝ��#�W�)QVF�;h�w1�~|X��>T�)� RU�	��J��F������hR�p���Y�/@l�,'f��Yt��a2+��#���tx�!��a+�`+�	qkq�x�K��ZZ�h����v��9r�1ҁ������!&т���crq9�%���.^�=���͉"�z:��x_�����6�(|�L�>�������["�zdv�͙�R�Ev�����k�5��x��4��B�
Gnq�H]>����HUH�iS�	�	�~:��Uu-��#s�j�����Y�;�D=�c�;% �o9h3�`��^�Kc��e�̵�g����'6>|m�А��[�*屝��Fa�ׁOD`|kٰT�}�)�eW�� %2Ƭ��cn&[��5[x�Bdճ���2E�	���`���4hܠ%+>�9��U���C>"�Ob ߼2���
�W�w�����Oq�%��1��u�Y��G�㙆����iJ��J��l:��0\c��#�x�������㧕mel�VhR��@��O����h58�V�rn\s�E�1�q��c�K�㘏v�MP��-��ԣ�W��l� @��FwxX2
4�h�ƍ��L�i�d����?�˞�V�K��!��`L�"�n�"�/��ِ�c�Z���!���=��\�Z־8Fkq�RM��?3@��O�����t�vm���4��Q�-�L�`b��Ʉ,���cg8�2���FfH)�	�'^���YT�8��_�r�ܨ�8ӵ�y0��2��Y�N�z�ܯ���+�b��~pƵj��g��� �$��n+�#/���Β|屍�-6`+?M�A!#���Q�\�����Ȳl���5��]с��o�ڽ�A/�*X R<%����3a��͖`I#�3�$��Kb�{}6C�(�h�YR��y�Z�ctPj~�����m�]s��	���j�_��a�k.Y�c��g*����^_��Ã^��a���pԔ��hc���Lm�1I$_������ɒS���8L�	�	8,^!�I������7�w���o��,��"oH׌���	�{��T�u�s��7��X+������+]1���@�9�fqx�A�(96�s�4ͥ��on�]�*c�f���0�h�UGs�*q}��:����'�f�P
PQ��Z6)�E5/$�tC��p�)(�{��<,cT�y���2��pyE?OT$% ����i HY���깳5/��I
��
�ݕ����Z����W��y֫���������`�hN[�5�N3~��. �'���x��i����D�>�iXZ���C�����u�M��"�������R߾lb���3��o����K��A+����g� ��Z?I|��zD�D��q�Џ�˲W[6SJ���7��!֙�HS��t����I�<���[r,e��f�E-����g/��x��Y�8��|~�~�t~K>�3zb3�^�8�X����!|PY��ޝ�~Ѣ����e�p3���J$�g���\/� ��*���Q��M�Eݟ5�fhj{�P�[��20��aq����@���K�	�
Kճ$+�4V[�p��SJ�U������n�fR��&;(:Δ7� ��*S�0<0�P�tѣUW�"V^+���\�J�́�P��Һ�&�M#���+�c̭�<�`ӑAM,�T��
�|�j���%��^�V��~X*�|������CQ�)��-;�
!�>���ID�(Gi���������v�گ�2?��e͜�jXEԑڌi�ݔ^W��u����j�m���6o�(�
lb �)jm� �YMf�ט����.�/���c�����L&y!��I���?�&[Ŋ����3��xG��v7�l�끒��Q����x&�3��V]�)�.��6�'���p��?-�AVR>uP��[:-�I�S+}��?q/�9�B#S#��$��vk��#���ƘX'�q�Ao�^	��7�gT?�h+%/������#X[ws��>��,A{��p�w��0�j8��o�l��dm�o�d�N3�ʰs��b�mwB�S2�7<7�ej҂nba]	i/̤*�#�R�G���~@.]6nù���tA��V�tʗlK0'�M�Z5���pT���c\l�`z0�(��]�y)e��O{잠��.&�--=�vnG��ש[c���dWכI9T�G��Mv�?�(Ϩ^�C�D���2[+
f��ߥ,�cZ�̿?�F�u�]����Ӝ�-���b*c<�l���"/�B�B0���Me���5���w>�Ѩ�$�NƘ"���J_�b�$��#!�~�c���b"�J�Z"�܁=�N��-Ǣ��Z�}S�}7^���b��H�(����j�GQ�tu*�m���TyA#n=|F��x>�V��F1'�I�R�L?�o�,Ro^/E���͖�"۩X/+6�~��aVAKA�fJ>,^�[*�Ԇ�T�ou��eA@4� �r��f��Ua,M�ӕ��;p�3�p`WF,���=P�������h���ո��]��eM�kM������R����KʐvP#A��1�z�ia�Y�����X����a��'��*Vx�Y��^'���޽�F����nOK��-��n�TT�/:�z�MY�HȄ�gR�+t�)M%���0��2��� ��G�/H4p��?T�K��F�p��E*���)�Gﲃ35'.ԫH�|3ݝh,=k���������*�@�rI�w��j�@&�B��u$�g�������+�����ľ���; �!1�QjK01��<l:��&A��M��d��ƒ��B�#�Ła9���t>��U}�Xy�AWp�ޅ�&��҂�פ"8-��-��皳vl��������޷�z[p��j����%Ӧ���0�!!�e�o�t�]�f���"vo�]�� _."����`]���^�b�9�p�L�0(���J�)q�`����`1Ĉ�h5�R��^d����6�b��� 5[���8�`�hQΈB�Y�9'х�1<����E�P������.#f��	dQ�{��5zs�Q�rI��+M��W+	
]l�T���:��"�q�|������3�3��rR|�4��ż�
z�1�0�����p�	}E�"1H�̆�j��Ϡf��R��XB����x�N�M�;j�qkH��.HDo��"B��b6�i��b�機���(��z+��բp� m��;%�����2���N�TN�vO��T���]89'�'L�<�!�|tC�V�zQ�G,!��.j�NA��7O�ż�@RRX��.ޭF�|�~��Ǉ� i]v�4xW&S.G��N$�HN���&�zq�|�۬7x��@�Q��<A�Q����^յ,��_�<�.�0~4�}A��\��QJc(�`a%ʂ��C0���h��p�/�eհ*���=K�@���v�ٝ���E!��ع��=�}M�Y R;2-�k3��G����XU����������{w�+�aj�.C7��/5~È�����N�r����_
θ4��N��)�o,c�E�*35�)UH�.�����K�7RY�U
�!���� ��GY��o��\(=~&+�U���Vm&��¿b��$LK"���)uY��0�(�����yuF�Ħ�wI1&�]���C���8�Ie�ĵa[������4�]r�Ǵ�&�:&iC!�}8�0��	չ���Z�:j���J�]��C��?���t�V�7Rj]%bY	����u��
�������V�1տ�7�V� v�?�0��ϸXL�V&��w���,�*R��>}X�wGv�z��C���+?v�2#�S&���i`/�[��WA�G^�  �r�6$�'�%��n1塁f�*�'�sT�*�u�!�S�+����N
X g�\G��7%��(�W31�� 6��n�J*"�/����ˎ���z7N
^�q��uͥ���������5a�j�E*�І��%�cա�������Y�J��NG����y�i&�3a�/��&d �8�����!��-Dl�^�X�ݮX$�"[U��y���c��i�Yѭ)�+-�2������q
�3Mu�b�q˴��~��k�yB�� ��P5��'�me��7���ވ�`޸��l\)b�qvr:6��݂�C?Pp*��?u�&����]�$���[K9�׳-#V^���.[�}Qr!�Mq-�v��Ϝ�WqDW�AT \(�X���
C�ea�n����O�"l�'­��K�����bi�O�s�g?l� �ǰ��5��%�Ę9����VlM�`s�G)%�O>dAs�U�Cl��3ِx+7��L����r�bήau���M���7���-:h
@σ�:G(\(wٶ
���\����Yjcέ|���%+5��D�h�?L*�{=L~_E�L����z�{�O����E�=M�:m����Ha��1�����:���kmU�5�>�d P�$c�Q�Ɯ��M/
.$�I��ě��y�5	��bh'�6��7���[����2�k-2?����B�!�y�k� +�����h�����J(J��$�h�w �Z/U���R����:vǦ l��6MEV� �t)��v�Uv���uB��ҷb
�[�v�Q��K��f̄B?������#�r�bv�{���6�1�[͐�����6N��?��iYqTۤ|C�#��b�� �n���&)0a=4M�p�y���˸���/�����N�F�5���3�o|��O �	��X�5�&�2��R��kmk�("4\��1 +���N)����)=��K혝<����@Rn ���{�]<&3�T@�=��h�9�zT)u`q��dy}n<H~{�+��/3�n��Y���&�ʾ؋������ġ��U��/����:X8t�1銥�b^K}=YN�30İ�;������C�j��\e�/8"�2P��K����^^��1���<�4��Unf�T+j�Mu��b�����d/��Je�`�qsΰH�%�L���Wb^��SQ76P K�n�wI�v����_|Q�*�i��K*�-�/!J��-|��˱��U����>(� G]b��x:p����eh�eνp��2��jfiv����>FI����7}�!�����+q�@}���!-P4ZtC�D�|�-f�)�{{B#�4p�;U�i��X�0���D1��UBb{l�����7��k H��@�'��eݸ�%��o��u���S�5e�_�S�\�}U�0~b��*�x� -n�e��!�����g>Ç'DI�}�K$$Ji+u�;a����.�>��֧RM����|ӊ��
�꣣�D��)���^���6q{�t��ٯ�U�x�ߔˉ�ц�	-�L��N\�s�8g�w�+��?��T��T�^J��Ký��wv���K�!	~��$N�j�z�	�b.�eR��s������7K�ϸ|r91y�9v>"�@��m��� v�C��2� �Á�ީ�0��טb7��,��GB��"��zѴ�^>�fϛ�(�؜T�>���E��um-!V���{�������Óvz/���8�tP��wZd�M�{RU�s ح�Dk6� H��\f���&��A�+p���������6�����y, �*jU#^���(�*?�A&�V�cE���?��W�I�<����>i�9����7�8a8#���wۗ��g،���j�U��Kr�	�u�[��#��b&o��(IS�yG��K��T���ǡUݤ�s�MCE#����jv�̡:-)Y)bC�X�DJ��|�TY�C}�����(z�p��W_L%|n�����)�G-��J\f�s�/hkЮ�R��;�)��v��2�Y��h�������l<=���F��M���۵��ӆ�o��d�5۷�\`�^���;����G���|cxE*-�%H�����������_9�ǎV��965f1_C@`*S��J	���S���Ed��c�P^��H���{N�|�q��_9Ʃ�͆�w��������ޤ"_A1�'
�ҘZ���1��a|��u�3�ク�"k���3C�ݗX4dK��H��o?K�;�)�&�=c��ϖ�jՔ�acJ�H��� ��;$޺e2�2�I+F���	�/6�ll�jMھǬð"kP���d�	��(���C�K���l8=Ǡ���L ��ɬ��v�Z.�i��sHq�C�\��J�o٢�x�����1���\�=���&�j�s)ST��Ϣ���3��=7p�L��&$i#���O�@�E�}�B�ƕ��� �� tr��C� �
�䷌�l��������D���-J�3/KXcD!!�LzI���_e���r�?6{��W��1H�5I�B�'J��	cr�]�Y 8�^�/^i!Z��qd�%�.��I���z��P?���MR�h�.�S{<�HhQ��ԕ>]���캗�v�Տd�>�B�ͧ���j���# ��k�$��-r�va�A�|/n��{iR��>ѫ_��n�k�gJ��P1���Y�6@�#��"�*	,�(��ؒm]�YĜ�D���_[�Zp�_�]�1v���Wvv?"�� �ug�-/jմ+�r=7�7��~���']^�b�������c���W0Xe+��<uSD�higqiX���Lj���Fj��îI����c�j�<�L0Z%$�5ٮN���{s�F�Mn�oH��+���qQ�1�yw,bu�A��ؽb[��A�"!
B� Z����l��>���,[3sj	�%9�T^��'_��L�h��.h�^��8��R�lpnW��S%(���fX��#�`�8�ʄ�l�u��n�ĉMN�i!�^q�K���hbAI\����h���V��.�����E`��H*�x\<?���?#�?�>�OpG����pc�ڃK\��&t��m-���ٮ�����G�������Mf&QD�����(��S�j�X8gV����j�#�*k2Bl�M�V��bY7+SV�x����ێZ(C�8��)-d��D콷�������J��C�cJ��y91 ��r������/���Z���%a���	f�ț��ߢ��gT��X��Y+�?�+�j��\�Cu;`��21��[���|�c!�1�f'��J(�"�wtU��F�٫�Į�`��4K|`lR�S�i
��	�_�~|�}��}�O&�YOV����IZH,���KB���5�`��d�x鄆;�1RN�"�y���Әɣ���>��uɆ��O��������hmH��S� Qp�`#�ˮ�Q8b@� y��b�DhJ��gm5��A�.�u�͋�t5\�lN��)�t�+�� F%^��@�-���>�����ĊF��X���9��}0K�4��dƖ�-�I��(<�u7���77t�'J�*�;7�ҹ]x@w�RSG5�P�0g��"W��x eDEN �؝Tgc���������[0-��
�YԒ	Zm��E�Y��7��u"�W�'	��QX����'N-O}(�fw�;���]>?��ε!\�rK�F�^������)�ٹ��hT�jN�.�qg�O����=�Ξ�%x����A;��1e���>=?cl�dn9� ���k��q�~��V��6�hap�|�@x�����SgT�<�	�\���"��E��V��{��o���=(�+�m/�j�'p��H@���j��=��AE�5�1X�w�����k��(~�r�"/�w���K8@�v& w���҅��h3��n?�F��d �:$�^���fF\�m� �fk)�?B���]�tX�$�JR:�/"]��?�P���:�ֱ|8��֤��˲;[���!/^d�c}qh��?Z�s�;��ݺP��~�O��~�6T��d�Q��%���i�����'Tq�3X�6�K����������*q�uC(ףs�d�qi�V���̞�8
�� ��'�?��*t��,�(�R_l�T��!ًJrW�+�5��� �����b#w`ի�e�[��P�P�w7�1�f7{_\��P��j����Qzf�,��B�qbU����Ӿ����2��]e'mA���X����-4��y�k}��q�v����.�F;yJnY�I�m�r!wW%.�I�;���ĝT�����N]�H���?T�vm�^�9��X��ǵ�������;;���������`h�	틟����QC�	x���?sv��/L^7�����WZ�S<��i���V��w}(�]N�d�-3a��p�x�U�#1�u|�:Ҳ�
�x�}i�7����Q�)�O�%F`�ah�KN��5�O�XC�R��iZ4�l�?��^]�>�fA�-tS�}�U;��>�ǂьJc"�m�D�ʇ���Q%�����!i�Ŝ�S߉��T���&�Ճ��bw�E;�2u:�PGP�[����oƙ����3eӊ�����͍e���
��E��?�����֤�02m g9J�~�A�Fc�,e-��A��"�u8>�+�v݆���h(�fh��������ӾvFg*ͮE[�ϐX]�?�g�\����D����A��7��'�� 2��S��Y�Pe-�"��<�w֘<4(1E�	ns����#��oa����ڔ$���+!�Q�2X+aU<{v��:ê� �kn���~9 ��� ��u�70=U���\zY&nB�S(<� �첺xv��S�&�JK��w�N�@�c@��Vq��*�֐ �«���Y����,�d"S@S�����)S�kZy�s�ڎh��N|���a��I�R.��Ss2�G{X�x>�BL��ԣ��jcl(ЩK�H��%�(p�`K�C��S���a60�v��Xk���P��7��>�K�B|���+�%�.����]�$��\J 2��r����v%X�8���A�'c����+w~Z�GY>���̷�Cu�)��s�����+��d	{��6��K�֑�k4#�<��+�.X&%@u`���n1�	y�b_ S���j��X�X�8ĽU6�)�����pV~�&Ҧq.��n�[�X�C=G���{���C2��Lb~�&^�(+�a�rĲ�D��a�yc4h]��dM�?F�=?l�;Ն���d��I��B����t-�{����=�}=#�W�⛱���|�M7��2����o\��>���ۃ����0f�˟�p���f���^�S�`���lU��:o-$��
kZ��Q�O>��XR'W�s����FI~��"ԪY�����}T������?t��ϝU7�q���N��zGz���_
��ȃ*E]��ɭ��C���.+u��-���
!p�0�n����OFz��#e�����Fůж V��	��.f�|oꐓ��P��vR�%ny��fq�^]?BF�_�ѭra�L��_������%�"��G?PK�nB0��~��↍��������	��	~2 ��r�T���l�d�S-���n��-�Y3{i�KW�b`O��Mʲ�;Sn�C�$o
��S�J���yf��m?7P�]�]�-��M��qT0���q�#�˜L2Qf��j�#j��ӽ�˪U�T��U�A.�����P�[�Z�\�+��X���iD^{]�6�?�	1�v�K��77���q�ݘ�d�?AX����)���F{N�*�.e�~��h��ٽ��H>Z��?��`|��>U���er�p/���^��B��B�}�DS�O�4�M�:����_�<�G��w��Փ�s	�{XW�,������"��VgwN�zL���ӧm�1W<��4���܂�.A��C���'�����ēÃ��2"�~�܀�m�$��w�I�I������ӣ��yB�3�jw�M�j�1�*����0��R�o��-��u�)�0=�r���s��T��s�n5��'S����L_�L�Uj�;�q��K�M�?�b4��7�"q�Њ`��ၜ(5���:AT��+xO/!A-�"?ZИcuW˭M.�{R:#��),��NTC1���ʃGv��w%�>��/����Цw�=�94Eh��`���R��Ҋ���L�*	�E�1�Ԅ!�r��iyd��y�i�"�Z]T�?��E3Fcލ���{���?���意$��S	w['g�-�DL�6h(�4��5�lV��O8+��}��d�e�����Y(F3�_d�=^��t�l�N�n���f�ݲ���&�d"7���m�<��J�)�0<g�
u;v��ژ��ʂ�q9#+�U�g��>T�cū������!pp uk��%0v6#7iT>=*��>�}�>Be�aGMB:��qj����z���M�fV����b�B��0��l^j�<�ln���4U��򀈫��؁����l-��o�f����=��#�6�𞦇B����Af��ܱ�:�<o���v 2č�{�k-�y�@����8e8�f�;�5��
aܿ�1jw�uq(ŋ_7Y��r�{-�^��ĉ2E��+ ��0D�d�4���bk���t�%S�2}�(s+��|Dg\p�ວ%�������MХ��I�7�ed����2�D�H2��D	��������	�/CT5(�(����O�I�G6��h��F�>�qx	D�#e����Qh�'����O�6��9�;��c��y�ɳ�+��]���H;��t�ZUـ�׎ۅ���"�����"�T��TY�I�|����=�#.]T
K�X ��iHH���p�ؑyJ�R��ll,��H��4^��Sv�'e)�}ӪJl�u%�uZ� �Uyĭ�%|7Rg��%	�p(]����Ƣ>�}�Sre��J����a�U�@7ꄂz˲g��J��Λ.q�S�a�2�'B/"�V@yc�<���JZoOf�k,��LNO�J���� �ɦs�� �,�����ǫ�ayތ�1�u���[����(�\��:���{9&"�V12�b�$�,����1HO S��>���"V��nb>pή�@��z�9���Ƈ�:���@�f�?tt� [���5��җd8�t@�a�0����=���&�U?lta�m/HHj=��l�m�0:Æ�];>?^�kӳSέ����3-@0���+U�g@�	ņ�'z������+h��@;��{$�>�ꕏ�׳L 1����|*�{�s����Z��` ��]g��etl�T��C�K�����E����	�1����Jӟ�>2ay_��9 =�O
yމ��-Z��7p�:R��ꦙԵ�ĥ����`e}˟t�cܣ�Ʌ�)����������� H����*�8ݛjK�Єl3����$�"P?K����n)9G���{d�s�፰�5��O�yrs��)��g��>
������`�Y��1Q]�L���\�*�ГT���WU�.v]|�M����jaLoǄ�|���},�1���R}��O��V?���$��{$j��P,`�Z뉧$���x�������5F�P�I_<q�� l��|��Z�V�c���jn�'�뷥ͥ%�3�쥧�����<�,+~����+Y��Ԉ��� ���|���1��4�z΃_�:�6BJ�,1�/b��d��)�2M���K� R"IkKZ#����Z��f�l�\Uj�*,�	_�}3kɱ	���I�Ք�J�A?Vڬ��!J=˓�6g
�dpDv3����\��ヴ�r�K��#^X3��q��9��(o$D�
�J��������ǔ�/t�\�O���O��V��p��̿��s����,<�Ml��
x�Ue�����z�l��_����ƞ$>w	Qmz�@��Bi]���Kp��ü�pA4x&(Z����n��?b�����7�}^G�%�ynV-���z(H��4��y��[��8F�[(Q���?��Ko�,�K��Q��)�A�� �D�� B ��C�P�ݡ5=��ѱcrݮ��z5	�|n�έx
۸c� �ʤ��4~DP�T|���_8��L6a�H#�jh���W�2��)�*IXc!l4�|��b3?��/Dif	m�"̡ݯO�:l^ŎHi����~f���e����b妚��o�/�T�]%h�����b���$G�A�6�q�`]!�3 �]�Ex�<� ������GdX�����9J�g�M�T�T��*
9�EQG?�up�`�5�
J�P�H!IGE�b�eX�@�x@3-Ϟ[#;�j훫#�[y�F��$ϛʪNI�l���7l�޷ԧLt�Z�ì��V��h�&�ȏ-�w�*��I�N��B�&���ƸD�^�&�s�bα�Pנ�i��{��jY 9��!~ʐPF��Ő���=��X�l��"U �����}V�1yΓ�E��A���w���Avm�u����g�Ij+�y\�k3���|�gA��\��'��'���ɣ;H��N����_��ةk ��I��r���V�CH��Ы����`���OD���ga-1�l-EG�U.�ދ�!�t�g}#��q��>Ua�|�n�@M>J_q*��ɸ�T:��2�KY:�(�2�W�Y���`f�0#BWw� �������/�:��q�����*m�OB`�5o��H��eI�KpEu�f��W�L����J�|&0X�pݶQ�-��i>R�UW�v�m`�93���2qG^��٨)��zē�}�/��"�8���,��I����9ޑ�w���˂b�3��� Ll�u�.����:t����R�yKNc��t���qZ�ݬ�fK	@	צ���r��	0p�p�����Y�L�(;q�"�N���
#�0����)J���ܪ�Od	A/ޗ��T�=�V�m�@�fc%�'j����C�wa��M7XE���sW��Ĳ^���,����J�V-�nY��\f�}�GU��VQ�nb��γ�@���u���l�S�K���܊��Ɨ+��_Y�n[ٗ#p&wm�KHN�CT��	��fՅ$�Zw�b�p�aW��VuS��lD<�8�����D/���Q�|�G;{�ٍd}�q'�c��{p�!���7.��Dǖ��ez�<(z�m�H%�����Fubb��t��%��"��+��̊����қ�;�ԿywQjP����59�|��x=���Ȋ��6g�z�.Z�Ǌ�$ia�Ҕk�<���	��\�ɱFu脬��&K�qʹnR;������dK0���į��&�˒�2a1\/0����|a��^����ڊ��ԏ���R��2�im�����͌қ���f���I�Ha\g�|t�ܿ
�ֿ�����FȃLUA[z�JS���=��3>�����l�֚e�=�ҁod�`�E](u>(��ۉ�mD3*�/;<�Ě��ˀ�e�xϦ�X���
>���;u�|��t�F�*�H9h_�j�@�"Lh��7C�&;4�4�x-��}O���,�J:��p�������ءx����v%?;�Ҵr�x�{m%���R5��͂wU�Օ=S��`�F��8��l��	0�Y�l�#C�߇�,�����������6�����@g����G_#��C>���z؊����b��(uǢ�J��0�=0��� �8���N����N�����N���r� � Yh��;J|C�1�Mh��Ș��}Z�F�v�
�Vy0u�0��F�V��5�N�of�)�a~+>���&0���H3O��C�t�,h3�w�#G|6��,�S�O.#�8����!���1�l�r��K���������Qk�Y�~���:����}��
x�Hq)q��^�]M�m�O���a%Qib���=�Fې~��z����L�E�w=l�+�~�P�9�0��X�3rGi�~Y=\������c�0��UhBF���Ƈdߑ��iy�{�1<��+��V�۪�q�s�>*>K�"@衃�Ja�ЬF��'���
X�������:9�:k�����#��smϝ	�צ��nSk�o#�V��-�/���qPo�#�S���v�n��?���鼞�NN���t�0lz����`��������ڮ�tA����k�����f�f�ֶQ�Ӷ��A`��+)���;v��F1�vU��`��)���R0Ĭ�zua�]=�p��7�Z���{n;R�cу�30��p���s�RE��tx,�������\JbU��b�t����x�`��wd'Խ���݂7'�����0��T(�6��
%�e��}�b�b�AM#�]}���0V�iDѩ�F�)u�U�����oc@�;�x�l$a�i
6q{�v\�����9�<*�n��d#��΍�F��:�����H�i�c%n x�8�㻵����&����Pk�Ǟv�.G��_�#F�>|s���	]JfA㶜
���d&�]�q�g�x�Dy�B�a.5���^�? དྷ��|Od�(8J?�{B �?'��՟�P4E�ced�P���3b�=��4>��)��3�NX���=�O5b��,��K�b�`��:MB��ҬN]V��^.�G��5�|,��#�#|���x	p^��ٙ��}E:;~�d�<rl0�k����5q���-���D�JeQ�ԳWl�����j�ɠ4����ޡ��SP�?�KR�����]���L���I�D�ə�9��Q�=�+�y�:&t0B�-�t�z�T�k�q�xe(�v��)$Y�Hѓ�Gg@�"���Q�ۙ��S���w��3�
i�'��(����{	�ʿ4�%
�Xч4/wtR��?�B����J��)\N�XCoo]ްi�&��B��)Ў��=�x����7�~��U=�M�y~��l��D���	T�Ĝ���'�_4T����B�O�a�qW��F�C[N~K�����hrQǆ^�KKXX�b��Ũʉ�	J�T,�����lӌ��mi��4<JP�c�v���fQqn�h�SGy�7�}@O�A��'`�cb n�f	\!���~"�)%������+Dt�ۊ_ݰ�z
�m�����V��G��3��ig#p���&�!���ڭ���ހ��- ��S� ��Iu���rr��eׄ������c�xVg�:Øl�A�27$:XƮ\Dx���%��~Ƞ��I��kZfGDA&�4��:҅WJb�L�{�g�U�����ka�`��U�$_׷yk��nVG��78x���LN���(�|���%�y[9U �	�����JӼSe����y�R�������vJXa�-�'�l2|�S��n	�����1��"e�2�8�wB:	*�
@��e_�*Z̎��?٬�b�E�>��fܾK1�?�QʜS���`D�CH�+y�
�r�<g�rO%k@�wB�Ɂ��1����b�D����)��n7�qʝ��>�;A�A~@5��kPBsE\��8ӺOI+8��0]pe��{p�`!���"���Z�@:��_�"�7�S�4�����~����à���r��Ƕ��ʬ�r�lϻ��s�> ����O}�c�?�G$���%LH�Z[�}\dH����úP)��%>�t�����Uٱ'�7���bJQK(�ͺ������X	�/І2٬���<��j,TD��S��3���\������2�¿4���C��Oy�h�9n�g�5���͍Ǻ�ts�^�έ4{�'殲 �9}	�N��e���P��E�f��B���lq��0'3W	����J��1e�ӗ���Ҫ����	��2U����T}N2:_�SH��k�����1l�� ,���� �_Q�	ǚ�f-(&vá6�	ߛ�h�Z4"�U���;�f�~�d�x��d)Pą'�c�0��F��O��P;L�����4ׯ2f�xs�^�4[���땧"��`�.\����E�+(��P&���C�h*퍩d�s�DO����1w��h��g@�t���ƭ����uVYu�m}��J��}�<���^#8�6��7:b?�!]��٫Iր�h�L�����R�
�œ��4rࡣQ��LO��A� }1�)��u#�ԓ��:^?dd�O�6��K��@�~���4Q���n���'io���=�p�"Y �Jj#����/�#44F���,FeN!C��K<P}��H`�K��H�7��z+���Q�nu��1�T=x
`'���1�S]�R+j��l�Q�	>�C��<�XT)KYr�;�����?!�,�Sw0�gf���j�q�&hj������!�B�4�_r:}���q^a4�BR�R�KA4��hv-PF�C��&�f��Q�,��X��]D����*�x���5�%�	�Ձes3�eT&b��c�W�,�v�6��^�±0M���������Rr41���D�C-�G��j�	&�>8K�V�C�Ə䬒?������H��Sw�ʏ��ӏX�]P���y"����" q��pS%{�4K�$�0�4��n���Mw%`>O�����'p�'��?	(�PYL���2Y������&]v���������$��!F��6n�_?M� �J� :�����7��_e֋��
o-թ)�������}��T�y/�L+���#U��[|��S�Oy~�(Xv�<�p�|'���6䟣��A����>���ޙ������A�f�W�!�z���.�+1͓����<��C�R��(`My&wpĘ�x���>��X6fK�oWG�%����O����{o��M�
i���K��9Vj�c>���%���P}̡��1�R��U�b�w�K��}�� w�n��O��y�G`���onu�=H2�F�`M1�6�i��	%ґ�.��0A�2]M�ؑև��x� ^�Zk@��M�J��ɨ ����!_;#�j��j����{�L+հ�w[��,+�t�kg�4̷K*�>d�k�-�$�In���r2ei4�4���j�@~����k�O7�u.F�N����_�6?g�pc�X�����V���R�ת��n���4-$�$z�U	��βB(�^���]:c��"��s�Eq��%�#Q�~dMғ��x�����1����Ĝ�G��iM�F"=��� h��~�iq�F���.I��l:X ����I�*-R;΃�Ij�h�%9�英q��R�=ъ?���Z@�	E�B��*�#`�$Av�Ev.��W�E�qNϑ�BJ�DeoU!�Q�.!���@�^�χ���<�kH�g���ɐ��Y7V<V�x5��#=�I��Dfj�f��C�О�Y�Y��*5���^/|@�bv�`l?�Wl<-I7,
���dH*��c��N�%��$�G`�ԇGv��y�`��.�Դ&;�h��SU-^\Y;	o%����t	�gk��]*���t����<�N�fe?+�0��y>��(k[NL����ޔ���:S�J󨦩s
�$���▹F��GzA�M,�*͑S�����J��3��Յࢿ�2K�7LwZ�W��n�d�ȷ��9�`A�	������p�&�d1:���V�k2' ��8���sFxf����!���j0��s��%[F�ۛ�]_�ǁp�4@�9�rD������&nG[:3�#H���CZK��7�>�r+����h5i�0�E�o�o={6��mb�@r�@y�6�҇����L�{�J�v��f"��O]Ը?l&n
ug|rsww�O�j�� �����v�/�����c�R*,�����B����0�A�Ԡux�0��u��L�R
9�	R�a�Q�͌���+[�F�Q6�rv�����!s��ʗ��-G���t	L��Z�泰L4U3�	Hnqa�4P)E�w��8*��+�����&�2���h�^*Ξ�!c�'�`fTl9��?%c��Ȼ���8|�`�r��+j ���Ō�2X�FL��S��2bbM��B�^������U(TҙX�x�ݽ�#`��m<-�kHe�8�ϲ|:���Y���Y�y�����v��|	�ҭ��17��Wf�R\nI����cǤ���R?�Rw��ix2���H�Q�|�Q��:%p r�S��
�@sͽ���o��w�F����E�a�Y�i��
L82B����(�e�bC���g�oc8��A�|4dMl�qmY��bE���S�틤Y7?dc�:��F��|���BIRޯ��;4*XܚB7��;�X�û��p�	�릸��qMQY$��݋xA[Jژ�B��h�fH�}����r��,*OF.�����Bp^ l�5�4HT�Y�� 6�i?dl�P�5O���y���?��_�Y��d��g��2Zj�5�^ ���Nݮ�'8����T�>��j����3�5���<�=�q4W�u�0⻟��R[%|*���؝��Z�="o���n�/K���	�U�����O�@}j��E�s^I��˶�2�í">u�ɲ�E�%᝵�2�B͎��]������׆F��M�ЈB��iY*Z�Od�SI�{��g@eI��^~Q����
wU���,�aƒ�:�	���(��o�
���2o꟬B��� ?AA��1Ō��Y9 eG��ܗ(<V���-L*]���2�F��0/��a�U��~�)[)�G0N�H�� ���S����9���w9�h a8*�}8GY�zFO����D��\�>���Q��-�Y�����G\��nKe-��R�V@���BD��8��d�a3[ڏN���1N�ܹ�m�<.���Qt�p4>�Tփ�w���g��~kD��^o
ɒ�3�lǾj�fOL�Y�0����M\+��߿zثT�߃�6N����U�gv�K3]�w}E_}�zt��F�Sz��C`E�;����+���jZ� &�ON��/���F~�0+ M���I2)���d��{0[���7�q�/�lUx?���▲�D�E���`pE� ,�#��"��!:��I\6�9d�z�e;2�8�D��~\�ɝd��h'[�.ے�<���φ��ʼvw�0���QBx��֭;�^{B�����u���8yd�4tu~� �g\��r/�Q��>L��m�3�St�t�=�"���b��_��hGS�-� ��@.7�4n:}����ڨ8�Sc�A���������G����	�T���9�g�w�-1*ʩS�Go?톏��;acL9"���N�`Ȃ�Pl�<�z��u�Ymy�y�.ކ�K�
�&@
�Ð��v����X��'�v �1�����ȫ�D�2$�.��:���'j���b勝K�+C��(���g-�Zz�K^��A&N�~a�wz��L���^Ҵ�<�)�uxhJCQ᳕����y��	����ZN���Hsu��r����@fkg�L�O2Ն!n�ngG���i��@џ�	#AGf�*ʎ�����Pff��� >{�ٽ ���&m[�c����&5p�(�N��]x�n��Z?O�����;ON�GRƏ������"�˙|uã�^�YW٩�5��O�ސYuF���il� �I9�|NLr���ly6Oz�(���L�Ar����!k�Y$��8�y���ӔÌM��*��#��gY��(�\��Ú�u]��S��Ԗ&g[�eT�'��]����Ŏ$su��ȩ5������%)2Ki�R�.�镆�f��0���3�(��c�֑�GGj�n�/VC���R�d�&Q''����s�L�	*-�v�����q�RfR���X�Yq��W� ��J.�3��V�ȚY@�q�۟�vF���f#fhwH�S�wVC\��q�ҫ�6ᜇ�qK�����c�U}Aɒ��?���w����Y �{�Q�Gb(4s<6��ށ�S+H��+���6�|����N����e�p��Z�,�݌��)�6s,��f�W擀V� ֔����E�=i�l�5
\�x���&C��	���f))2~*K�:�_���M}� �rIq�XAr�Z��/�����1/��P�x��F7N���z⁘̶�~�%14tY�Q��j�g}�BQ���x�B�r��O�Z�2�J5Joa��4�J�ld� �~��̚8����l�&�"]�2枟���R��c�(�@���$3n��X%l�t�<8�,X&r�P���{&H�Z�ɁDyv�x�LxπBOB��~X����Y��.��`��sx� �5F���=X�!��=O���*����4��፱�P����th�@j!�G�<wW{������/��g�+�Z�aT����d�]����%4nn(����@m�	�������1��CHH� F��:��2qL�ք"x��4��4+��2TE;umd($���Wb�5�[�ʞ�ˢys�/��O�堯ÿ����ʁ�G�y��a9�bK�Xj������1���U:�ʩ"��B��)�Ek�%� �T�	��a��QƧ"(��Q� ��������mg��d� ��a�-��>��5ৡ�sd@Y�����h��,-!�wp`�`,3�?�Z,��*I���%�,���t�S ��ql!L�hP!CNg���c��Ԍ[�z�)�iM�Z)�>�"�:�>�|���*�]&G>�qc�X��4A��u~�������@~�F�쎫t!���
�m)�*���"l�
�/%Ȇ�<���f
�|�%<Z��z�ZT��B��ǡ�f��1���~��0˰���J�F�����Ϻ|p�u�I2PJ`�}�R�=���<��D����[O�?h��"��4R�Dbm`�0��ˠ-׵o��Ì�ªPF�x�Dj�������7�������~<��2=��3�a��	�,{gv���!������,��;1rȉ���̞�vbe�7\&�#[
p	�H��Y����b��ʅ��<	"@��(@b��(W�]?�.�sZ����ą9IՑLAz�W6����za=ہ�+�X3��lޟ�� ��[�S!�4�fh+��5��1���\��'ҡ���.Nn�(�n���S���œ|�C�����֐�Ax����S��A�7�����P'(�P ��H8��e���TŘ�<|g��l W�R�X���`�
�'����W$9Rv�yU���A���~瓞%2ޅ������z��F��w�&eA%S��b`|�<�������*!�22��:�P�͘�Y�z0o��<0rc��Z��� N@��8B,�v%���8�ch��Xj��ɶ,N��yvx@?��5�F�����E(b����3�����p�Q�D�"U�pD�t	���&b�,QP?��>:���z�J�~2C�h�`�g�`9K�`0E�;
$i��?��$��K8)�x =�J	>*�;è�t� �fcP��?��^%w�>!�%˗H�g2w��Fs�weL�= ,���;vrmGOG�+�|i$�?2i��5l��@@����Mi�u��<O�ksj��.�5�v�w�6X"��~!c��h�yb�F=͢�"���a��yt��X��y3���Ԅ�q���[r���zę�;�F�QII��. /�m[��$ �8��ia��0s�[,���vu{�7��}F����W������5��.ׄr���g��E)#y}�!��<%�Z����;�%~@`�y��+ɹ�ha�h 
3��R����}ط�h$,YZL�T���^��ޘ�p��,��Ԅb�d�rm�B1y�����r��K��*���h��K���2�Q��d5	! �&v��aϢ��O �Bӄ��=P���e����|���6��162��x;�~sta	%ccŶ)HJOOA�6��Ox�Ffh��Cj���xqb��+�4��:Sʨ�� lj��˘aZr���t��?(�$&#M�@��7�r٭�3���̟��y,���s�����h@��b��I^{w�${��+%$�T��l��
SuK
"e�~��\V�NAS�:c�x,�)"N����������P<�Yu%�ɨṠŅ?��*uls+�����'d�J�N_|ͰVxJ�p��S?ˤ��a����ZҺ�����(�8&�hEe	���yC�t������Un�3.�	<~Y�=X��<����<k���\�D�`�^U-9�>eN:pRi�-�}Q��%��h*�Y�q�W�D�у�JT�?x�*b��_η�}�!ƚ,S�h^����P,Kx�r��������A�3�T<|��"�r�ڢT����;�G#<ނV��f\��>���
��N5k'���&k�b8�ʾ������������eWn��Q[���]�N}���ҏ]��ir'G$��G캣/�]�@��&NԜS����h+�?-��ق?�hf�>Ru"ٷ�З��E�k���o��v��*����'uԣ#����C���L����L�5��CbO�xҽ��9.�Q��dW�qct����:.����)��t�M (�6��W�;��գ֞��$C�r6@`����N���E�H�F�����cO`8��O��*��A�BgG�ie}F,V�yj��D�,���v�����}Jm�y�t@E����?'�w�=_QY�[� �j79W�e�S�uy�?2_�%jq����1a��;D3_�.�̭hr�U�E�J\�얷�8�r���~Y��F�Q����Dښ��"��{-qwT񥢑��Y�g��n���.�pJ��Q�m�Y�i�sU�Z	�͙dS���j�����lz(�y���l+��|�ݷ��y��>�V��`�?��(�7\rf}����}8j�;�:���}���W���\"Z��Ɏ�s���)�N���~~5mS25�ܮ���:��y�������u���*�go��kD�[�'؆�8M�>�X���W����t��.�ӟj%q�h��h�GH�����	��^�B����(Lm�z�J���shǫ��]q��߹��=�I�=��Z�'�
���YIJ�l�f��2Q�U�:�دz00�z#M���,�ͭ�WNCQ�n��a�G)������0.�LT��Sa4�����e��2�``H���}:���~�k��A������k$�JXk����ugCw̻��5�:ok#X���=�\7/#�����Ftf.��`�i5�N6n����Ѕ�*�y��DI��K �Tō<(A&/�e�f�R�)#Wu��M]H��]X\�6�2w,��E;.�˰4-��{Pn�:�¾bY�3d��~eH���\d<���,������Se���*��p	��(�B�0�dE�4���SJ��7��l��	��-k��d?�n���2�\�^�.�}(cg6���eC��j��7<�!�V���q�.�T�hg[�F}q/����8�FV�9hs�D�������X�G����Q�O�� k��C��G璬��=���/��n�c�v�i����$O ^����joߐbD���;�s��b���G�m �\.k{��W~&?��M����{���\�i�ťb:�4��Eb�i��v�cIH�J�y<����o�H�y/y)�|�m*���(ܖ�G��E}�}�g%�\�t��P~\9�TIl�]�L�B�}{.�x�&��I��v�u�ǽob2����5}���f����*���K\�C�����#�v�i<�����.&<���m�'�����F�Sf/m﷼I�*ѦkOV�W���x+�j�B+�'��(���v�h��e��lm��� �U�l���,�� )�3�-s*`E��\��i�H�m�h�_yJ�VA���T�m P)[�o���4r
U�@&p\�fܥ�/�`� ���������N�����zg��n�<PD��s���A�r!�9�~!}�o+Q����+�UT�
#�1Ot����+�T�0�̡��ӣ����~��qor�Q�T������1#Dy���F�U}��b\�E��˴��0�!v�BB�z�<Շ��.U0U��	�4��@���vBtf�/�weg�P���F�i�0:�Y����c�C��� !�Dwrl��aX���6\�j"a�5z<=��ra.���Z�jH�jN�X�#�U�bie�%`����%�rz��0��"6&���<}�(��'���ī�i� f�����L�D�E{ě9��8$|��%V(0�_	����X̐�4d@�fP9s&_6�.���F�w��;#�\ﭣ��aOJCſ��������O���Y��[���������:�҃CƑ�0`��g��[����xy���A5Fȣq��.��� �J�u�
D��M�� 0���(�H�[�g�l����ϒ�u-���((��[�ҏ���-&V>�@�s��!�"¨yT:��\7�Z�i�&H��"�Ε�V��K�Œ8�;U�}��D�J_�DP4f���~��z��@�B�N�*��;(��M�g��+�(�f�uO4�^��[�a����0�Y*���,O�]�Ĺ/O�2Tv��8����	du.�4��r������U[߯��W���ڮ0���Ot�O5�������W��YM�kč�����as!��1�Z�&}��n��+��k��E�	6��p[�d���D����IE�<�&�����~��B	���(��f�:�L�U)����5�v�O�6�Ħ�tJ�Z��IƧ�~6f��%"�
���o����V�1�T��Q܂P�@��,�9�t�J5���$�]l��yvh�
	uF\!�J�Z�����4�]���&ث�P���CJȌN|�Ȥ��acg��>53���W�!��s�=�e���p�j�[DNa��̴"���'��^��	,��*k*�X��$�^x�攔D���j{:�xؚB�#��X���G禦bh{�%�?�м��#(�:��ڳp�M�ҙN��1s=A�#�qi5\~￸h=��)V?�i��a�Mu��QN��
�x�U�׊�.��ǹ�D{�\�̀���򞤥�h����J����e%��l1�G��m��~R^�]g��+���rSj��d�c�2��. #ׯ(P�M4�X=�j���Tc�̛*������^3���Q�˵�]>ڿ�'���a%2*�*�C�D͍#�~h������ͧ�Y�ك4sj���L`eKG��0����\��S>�GWB��U��c2tM��{�	�B�x��I��i����_K� �5�����4�N�Ro��Y��Y�A�~�����ɏ��^��q�p�1~���i���o���:���l����@1��xR���b��*e8�����m��C�O #:���$�$�L�n�t�o���,�VKN��9m�ꫛe{m1��9���&Z�T~k ζ��-,w��ah��=�t4��e�}o3���ϧ��`��J�c�����D��hkO�hVa�瑦fV��@B����N��t�)ro?t�1X}�+,?M$t�����#g��z),5ɩ�C3?I�]=V�/0�J&nkTΟw�c,��d��~�U��%Z�����	'DV��Z�!�Wμ��`��<!�.5��jH�i����04�,;E���ۿGm�Ѽ�d[I�+�37U��S)6.i��O�K*�]f�]<����z4�C Hb5e8n�es�J?�Fnj;ЇxC�÷57�٘3V�W�o@]i�@�U�	��`�����U=�F�E1d@!�!���^x�5�]�����C���,^�T��ڛ�Cx,Y��5��S���c�@�K��xg��QY��\O����)I��$��ت�aV�0�}9d�y�+6���B�^��z�*ڼ@f������"�˵vg�Z�.���
���φ�h�&p�vn�b�f�n�>~�2w&��و5��]�",��~Jrrǻ�R��#�����Ȇ&M1`h�
��QIj�d�Ki�,�[Z᎜<���������6����D��x^E#��[<�xW�h���tw�7�Ċ�`��x@��K�i0���)���G��OD���F�뛻�&����4���}&X	�+�*MF�+~�R!����YJ�-Ȧ�Ɗ��I/V��4��R��G�g���f7��̡7/��r���
�;��c�1?���<��;0�(H}�|��H�1�i	��(7�#x#K�٭6��9��2�/��Z_n�(�8��)���u�����΋�S{��h�>��H&B��D~g��C�q�ٖ��	�B�*�}������J优�	Ħ��T��������r��� I�-��?ɶ_]Be�' $�@F(K����+Eí���憿
��B��s�1���{`��0�������f�EC!S�=�"�<U��}��glx��d<m�������0�(HH��3�sF���s�)Gy�!!�����V�-L�η�E���b�x��)Ⱥ������<�iq>T�P]���b$9{Q�|h�xo����Ʋ��c{|H���Y2��˷����j:*
�	mDvzI��2�c|��E�ƌ�$���plG�l�~l�2�0�"M�sٖY���g΅�)�u�_�V��&�x��������L�����}�';bwp4R�E#��d^M� �T>2���J�H_ysM+`='��:h|(�~V��AЭ�=?���r����O�J(�����������~��{+;9�%���{'�~5�7E��,���|��������)n�
=U�Iz[2��C�}��R�z-7,��X ��g����vDS׻��a��݆v@���K�W*Q&Ī�1�)�F�i)d�m��jI��~��#��Y����p�-�-k��m��7!<�C�w�$: .`�;_��ê�QB<�p�)r���6Gܢ#�`�#��������L~Y)��=���mN>,јK����-lE������[��	�(r���� _�[u*m���  ��b�_�AK�����_���*!:�j�����6},��({Zj�9���#V�W�{�����0��Nt�(w��J{���_j)�E�<�\��}�8���8��n�7*,C�����h�|��N�z\�e��~��.�c�/bۑD��A���WU���⭊ŕ/��C@f�ڣ;SH]�<�>$�Bש��b�Qg�������j�\��N�<�E�ʏ;l��'~)%ڧw$������3�w�ENJ��V6U_u_!��ܜ�ѩd�b�Q�C�Ry��6��	i�"�8���,^p���9��E]������C[Mf3\�C �\��)ϙ*��K?��s@�w(��^� -U�~K��}s�B�P�78.��Q��?#����\f*-),q�mR3(~�s�ib0����4�>�`%��F}�����Ǯ>v�2�&^�h��S���6\	�G������l����a�y��>���݂�{Z�X��o�=٭J��9}.K�́Oq\�ySs�8?��O74���ɧ疰�ۛ�u�t Q��/y���a��}b;J��H��[:����l����U�f��fӊ�}ӈd��CtPz2��u�>�u�p�o�,������M*��E�^��Ёi�!i�:^䳟���j��K��'*b\G�\>���d7�Pw�<����w�}�k��r��G� ��� �i6�հ>u��v̽�wVN�[:�b?�Ƞ�����o��|%6*=3T�uK;��'8#E�o\6�s{,į��d���`Nv%��������ב*��qE������O��͢ϳ�8M<g�4��j�8uf��:)��S�3ޘ���ι�?G���&����dZm��@���A�����>������}'�l���ٱ��ͳ��Z?�AEё�'}����Rm��`o�v	-D�^�j�=�ld1W��$<�8��9RK��|ÿ���02,r8��:=��MƞM�Pҵ��Ƥ=�j�F��e_țQ�U�h�&�PPp�^"����vF��-�W�����������Y���Ǝ#L󑪮����G`J�}u�H_ QP[EL��i��y�ѻ\e���:`��r :7N�X��C�Y$�w-�$s7�TKBS�=e͚�-�>e��7�w�����wM-����<UxɎ�l�-zV`>@������v���1%_j��Q���DL1����
�OɧbOB*7��ku������-��k�)���6$]f����R�nu�@Uܶ5�r$/��`Uң�¥z����#�^K1B��ja���"s�516i�G�KU���� �sN��#rޯ�zC�wH��H>>7�oj�'k�ʉ9����
}��!3�5CS�w�$�u����$I���Y��ou+*��S��Q&���~��u����`|>�n��*~&��J�[A*�P]��5��ёņ_Is�S�!����=n!���Ok$krQg��6���y�V�F~��4�Jϴ)��Z�P�P�������-�d���>�����?|�DM�t��0hv\� `ޔ�gsc�F���A-�i$o����t�]�t���j}g�G!z!�,�9Q�K�Q�m �^� bT$�e8m��&0�+H�4��r�EN��q忬�[E`\w�����$~Uk�����c&�Ma~�1&]V,vS Jc���3��V*;���6�m�Ԍ�Էv�5�AbCs�����	���c��Δ�["���uMSY^���n����c�Aur��|����8M��Ð�@F�''I�p���\�s

����;Y'O0C�K5&N�y�;Diz2-�e��pW����|��e6}�����W���ލn�x���{���I?�O>���D���5�*6Zs+�(6����(�?'�m��L}�v�*��O�1�2����ڔl�+7���9 [~S�'GH�!g
	��W@谬�ej�}NY�XG��ɏ��y���#�c�
�9�F���]zM��w�:���t����4V!��Ht�y,'y�<9U����"Q����2|����+ӗS6�ŉ��f�k^.���t�$8�/3<�]��e�z�� �r���`�&0u�v��\Bg�U�á��}~^�6I��I����[��a'>�Z��SK!����</�l��=�{I�y��q�_=;���c��F�q6N�̋��}+�m�iC��X1A�_�-7��㚮w�E;l��KK�B!1��^�&���]�b3� :��8���9�,D�faJ�U����������F�Zm$x}�V{�Y�#��/�/���yK5Iʣ
,��Jr�zJjm�mL���_�'��qv�:�p�S�t�m��ۙn�w��:at�Q+����L����b͙0ѐ�R��ϊ��ջ��c����/e���jK-"Ҏ0~�X�1(�o�����c��	ݕlA��o�	��������䢬	�i�V��l3D��nD>UMS5&��6�Lº�m�m���D��63�k$��!������55���B[[#Ve�(J���/W#OL�Z�}`����ξ(�Z2����5���R�����4�M�@K���#�9��WըN�5D�%D�h#���r�7-�0���OP���9_߰�ԋ�*skG��ل�#�\���j,�%��L�|r�d����Od��b�?��j��Ǐ1}A���.�P��r��{0��~&���]U��|3q?o�Z�"�I���*o��d�I6�� %�R�E���sȑ/l�y�O��%L�n�5F�L���4�w�ń�=���ٛ{� ������VP��h��Y��Γ%��]}R:�[�ӂ�RuK�u�/P�h����đ�h��і��J�v%��T:0�tB-�TR�
23��,1�5{	�i�׃8hf����j{�����/Qu�Zg�����h:��1��H�GoW�71�^����>A=���dt�O�.9�m���<�+M��Q�r�_ W��X��aK�ݧV ��UU/hI�����.E!XHۂJ��6n��
�����?�e1>_ĩ��}��)Dw��t)�l�q}*HS���r�T��SK�|�D�ck=����y�++������Ԅ�*�tpM)C�`�H}O� ��=�?�\A_2�v�]`�*{�V�m�T��� �4pr��/���f�ǝQ�Q]-D�Yz���/����ZoQ���=�<�b8�h��ܳg	�b�o�w�$
m�SX�!%Җc��ʾrk�"�b�,��D�b���<M��T��/n�k6�q�dfJ��74Sٌ��˪T�Ԓ��h�0&�����w*��Ǻ6/�r�����n�Ēʋ��Ls϶��-��=��.W�e	ƚ������}y�;�d��vRY������ ��! ���3d��^����0�d���2v�F��部�T��Z3�6��[[S�M;F�X�o���NK��6G�ca����kWU�0��WY��b�ƛ����q�:�&����s6]�
�Q��6�|i"��+��|~_0�L�-�r�7�%uQ�:�䲺˓E(��d�~�o�<�钂�-ibeM�0�#�Mk{]p��?��V~1PB�9�.Aݬ,�1s&S;��A�*}��	��]���sѡ0��
��0���г��NL7��@ks9:�@�
$�$�P��)a��. NR��
�����`�"H^ݪ~z�s��IS0���(˦�R"f5)�IAoxWV�a=놨ۡ�[�z�������I�hВ�:_��!��nn'����fd,�`9ٰj��>ړ2[�e�L{U�+U���g�r|f/��jg\��-}vf���tg1m��/�V�{�ſ��I8+Bd�a��3U }��G?ۆ�����R�8���n�T3i�Ư�����d��;��?�q� źձb�`9�+0�Z��UpZy�r�:��K�+�I���1^��?�!�Ǳ-JH�x.���.�ہ&GC���g�n�F_;mb=y-��-h������~�~������x����7;�<���M��#Da% �XCq��I̍yI&��!�lQ^=����+O�����ޔ~�yj������3��b����:�(Tk
�24�z6���f*!غ���K��d R�Hmy5a��!g�ʕ��3��'}( �
h�8�&b=��P�"NM�,�_`�RX�ݼ� �/��H�R�]"t�}�QԤ����C����¢��$g�(�G�ч�H ʇt@{���P`qD�tĐ���4�?����� �E����>�i�b(��4�A`�Pa��H�H�4�@�}�Y�` ��;�4_�y�7�B��⤄�˃v�ϱ�ͷ���7����mc���(-��5rGE4�9�%�s'n�<��"d���f�"�.�.�)��ͣ��2�N�7��L���UN�ה���cb؂iY=[� ���n��`��,�M�aȪ����X-,�?�2О��Oa �G�{ǿ�>�ZF�<b9	���f9a�.��,'����L���	��
u� ��[��͓���@z#�k𹒥�ђ��k���|l� ~�� Z#L�r1_a4{DZ/��+c9t
^-��4���E�����0�*%�r�ŨЗ��UO�@GlE�'"�S,9ڷn�x��`A�"��RD��$���4D�d"�@8�u�7Q\��[	�h��G��N#��N�5"��R��?�������_XJ��#U���o�x�h����~��Kq�&���,*.�"�SC�8�x��z����8���:oM#��c�-'�{��4�䥚|Hq�=΃���y��1�[��s�q������w>`��:L��ڤ�8Ԋ�դ��탽�>�6�<K�P�n�;�H�����R�LY���*�-*<��j/�$80g��<��ϳ��������64�b'��q 5��Uo]|~k���([؛F���&�ZI���f�D�Έk�L
t5���cm���o;EI��N4q�>ܢ\XX鿘��г�G����9�����2�Gm���$��KV�,�z�En=n�/��\��a�"i`X�^s�	D�2t��K�ö�ҋ����Ⱥ��bD���՝p:�w�a3���ƹ�$�6&�����J��ՁO*�}�h�#����߹�5�e�)H�3����a��z�8�=��J�wS�U��ٺ�����J�ME���{>f�����_z��kƽ#3(��}��T�?#�<����[� 5�Fs����G��xap���]�%*]A��M�f7{�����^����ԉ�h\�o�=��F}��g���S<��5�S��C��*u��6�n�]]�V<^Mv"��E��Rr�Za��~e��ܦ�ސ�az��Ŀ&���Oo򐝵��iF��������R$\��\@�]շ�4d��}�DB�l9��S��7���]���B\��< Sv!�n�.�1L,5�:��e�H,�j\�ŚZ�!f�Ʃ��ɭ^�WnO|�`��#svM�J�M����Nfߣh+T�&�w����;�G���	�4�R����=�:��6�FX�Os��RԞ�kΧj�ƹf�r��I�I[I2�4��vjB9��G��y��Լ�+j�G&C �d�$t'��=8�"=c[�yZF�K�;/�����}�4�<ٯ���#�? ���U��jχ�A+���@����-�q��*���S��(�s'87���Z�]��( ܩq1��<����B�Bo�]�-ѣd!׊.rLxj�]��a��!YE��	x|W�£[DS�*� ��C�� �D%`�
wIsv���d���W�d����u��ybO�`�e�=|�k(����R�Eg$9x3��w
�Go�e(�L�c�ȍN�֚�_�W!��n5���<��<vq����U���	���~��B�]"h��|%�/hl��E��j�L�|v��0���z����O�Ƴ�ٴ��`*��Vװ���l�
��k���o�.�4+����s��,l_�9P���ǃ�1���:��D�?w��J�7D]}H�b᨞�Sj�t��.����*��i�p�V��2%���C\���!��+)���0  ��_�>�O��]^�za'�H%6ie�y�qrŪ>=B ӵD8�*F�"��M��# �Kr��Qfgt7b�0���kg�q�+���ui�L2�AN}g2��B�M1���A��m6���f�'���u)��kBr-�����Ht-?
��\20���C�3:���<|��/��D��OUW R_m�� t������F~D��#�)e:>c�?��N�f	������=����Ac�������"����픞��`�4��(���ɦ���-��h%/�H�j��LMX�٪/M��r�����Sį�Z2�Bb�=;^��ɺP�K#:�/j����7��Iu�ݶ]� xQ"t�	�]���Q�#�/�u�D�'�9�� g*F ���k�W�;:Ԉ�g���uuU��W>�)��n�]�-kU��� o��G�*�Z
�<�Ν���ѕ)#n�UxA�<���&��Y�H(�tkX�C�~�3�/fm8$'l���r{�zӚ�}%�!���
Y��DQ.�����JD��A��j��lb��+_	�x���h<Ѵ�A�9-Ɨk��!7�Ѷ�h�#��	� �n�t9E_��?���7�ٚrM�ޘ�*F:��?z�������1	���8��F�CR-ڵk�$IxS�޸��`��L�9�f�j俢{�Y�h�J�JM��`^�ȩ�%e�+��9]�;	ѷu�i=�Y��)�n�L��NzeJP����/ed
~2-�d������9YM��ч2������5��\�#�M����Lπ��E+9&�wU�Q�w��S��z��R/�f@�q�`� ��o8�@��])k�h쥨'�O���?s�Р#2�YD�@��0�j���Si|JܱO� ��N�C�R]�߮�� ��R�3m��?�������7eh���@���am�ʲm�/�R�g��W�3��;��[��(�H�����.û�t`sp;:�+j肐Pw�c����̂�E�85�d�*fd�R�u��@�c+E]Cɵ�{�&�A�F��k/g-�6!��[�X��}cwa�G���N��%��	��1J��� �}���ٚ�����=�ԁ��L^"1U`(����0�����5�&fAj��8��I�2��5g�G�1�S���IGJ���9��7}�|�O�$g���*j�q�s�8�ߴ���N�;e䵷ݻ�٠��d����'[Ds(oѼ�ކ��U�VC�E:��v)��؀^���[ӹEy�� �$��}+�d��̍�
AeH����h��͑*�oCd����ƻR���1	�)C�z�oz��/�Δ�:[�L�x9��� �!�΢O����}</_���i�'�"�q#UZi
������h�����*��7�О�Ga������u����N�������p]��[�� :���K��H�#���ժ9�|b��~�,;���ѣ�~W-�۞�.�k>�HL���)~�Z��$9�=u`3tt��WE&��Zpm���'���[��|�4���rm�*!ǀ#��
�+*�d�gr.�b@��DH<��!8#�qw�0����Zޠ_�h���d�T�}s���S-i�bcԖfr��C��v$=�s
�pnt�&U��s��&�_�ָ7�x��'Cl[p�*���W�>�i�lW�V���(�^�lI3ѳy��A;S�0��>�89��$�	}w�<��Z�H�g������`U�_�P� ���P�5_��r;͠�F�]F)�sT��������r�6�m��P�S���~q�>�aϗ���3�؝��9F�w��i	�c+����v���/�z���%$�dAXcrv�h��b��Ș$�c�7�Ѡ���vns	y�Y49�{��o㫹���2_�8hۿ��;焜RJ�K�8ʮ��Yj�l��h�Q�z��P�W%��>�j�bPc:Uk��U�P����fYx���%t����W&A�3s��+jE���0���
4����F�HQ�PخD:�ǦW1TVaZ�R1@� �d��H� h�>���E�j��uQ�����$f�Ք����5t7JaA�_�c��v=&5���s��-mF�,H�;3��h0Ewӑ�"S��,R6
���P9U{��.�bY_Ȭ��RV�M�s$;�h��'#%e�r�������T�;�ZKϤ�>�BM��vV1���ٱ����K��їO�zX�e�+@�4D��i�E/6,��9��>fplť&F�BA���O49�z����g2��q.�yT,�<�*��� 7w	�m��@����koɗ�J�`�+��H����Qø�n�R7T�V&���������5����=>_hV�ìQ�"�N����P>hNJ��u�z��x���%�<�Y��b�˂.Ĵ+Xad|P�ϐ� ���y]�z�sls�Im�`��s\a$�5�i��x���"">�Տ��<�,�m��]0?��1��'I���G��(���h'�'8�t:��`2$�#@�&���=��1#g���1�F�d�g���,.�{���m̕�}}�d��m.�o�2J=J��o';}�9D@6�	
Z|}��#��'a�8���/�ؕN=��n?�q:�܍��H�l"����Üg��ï������l�&����+�]MԨ?��C�&3���i��4�1�{�2a�1/7<T��}e��Y'���ī����
<��������c�	��ҟ���vf5���T^�,(�U>���ވ����y]#�3E%P#b�R��[�����v��nk�I����!��/^���[y3�.r������r<.*T����T.#W�ّ"����_��ێ����c���>[���5��D��wy>�������+P�9� ��wۃ!��f.ꝥH�ېa����$�֯�EB���F#�t�gSO	�������L��p����UƝk`ܢ����0�b��z��@�J�RN%��>����߯l�8�"���6��CY��j�Rͦ	�����}�~[�C0�v]�!& ��ž�J�܈'~���8����0��1�Q쓛}K�dP���E�:f��e���rٳG�T��?�N��8
B�K�D�FYpb��J̾z��TN�l������:�+D�b�A1�q�z��D�����`�h��o�;�@Y�՞'�_Xᔲ�*?\o��98hѧ��T❇D�BT.�YLP���K�"Cl���g})'7"NQ�?�ԥ�|.����|n{�8�}]������C�V�w*w��ի]|L�0�8�-�YT�H)D�`Ƿh��R�0�v7��YK4RX��d��Uj���ӊ'�x�MQ�p�xw��s�[�	\�G��:�ˊـ�zɉ�i�
ow�<'�+Ug1̣�x9<4K/1V�T��ii�ha,�t����ǵIaI]�����n�r�"�m���0���*A��|P���[_�:��'�+R�!9,Pig��^`�� �i��eB�A�C󢍣��k�}xi.2��\�p���@�Z�w�jLy�ڛ��M��4������qv�����{�a�o<�.�Y-��I/�؈$~�� ��@��խv�k��"����+1��s�̸���ŚǎN� �(��W1�a�W
ݧ�
�9�]B-�c����w�֬%�`Uim�mq3%F��c�<Ș��Ԟ{�p$�3�K���=	���Xa��X������W���1c��3K���~Ձ��?Bcr�������;� ���S�Wܗ�Rf0�]���r��jTR1%�\1�����V��
��x}r����|�E#_m\�:��ծ��"R�b�C��^���*u$�,��%KGk�6�f��>C���_5UR,��>�;��0閫e�P6�3=f��ϔ�յEс�x��К�B�����wW�!K3T+&�Y9�L�E���)$�ךW�¥�o��9�V76 K�$��x/��Gްv���p�A�e�+@V�j o-�6�;������<���R�������Z��"R�Y!��q]�Lx*��񸭦[�w���Oh<8h'�!���V�8_96hmI]���,����Vt���j�( \��U�J\��Ј�3���x�x�L������}��=���YƐ�k�uV��yA�v/U�>��*�Tm.�WNrW����T���������u5����/����lLro5�Aί��bq]K���S� p�*N|"�l��t���V��P�=���pUd��ǴM	_�,3r0�8�R'���P�ʁ&A��z&g?�g2�S(~�U��� s>O8�1���ۣ6+���H�������1���|���9�P��t"�o��-������5`��{M��R���ˡ�hY�<���d�`�H���e�b`fe�Պ�w/��\��N?�N
�۹'d�S�V����k��~���x�o�q����wW~��������Z1_P��A��f+��z�S��O�t���u����n�ϭKcٖ�w\��"�{f���A0���w�B�<N��^�#	7c��HԾ0o��
rp���j�Ͳ9d�g䍈$����q8����9��M�[��:]Zܿ�P	u�aU	��z��Ӳ;Mb�3�}�%����,Y�fQ9���>ۀ�@T��H���	"Y���������7X�����W���T�.�"�ǔdN���&�*I�;��_oK�% 2T@�"ND�>n����I��
¥Db�߅|����`Uc@�8D+ħ�=V{�[b?�%Go�H�����^����B^u-[�c�N���?��̀�����8����<� ��h<�F�ҧB�џ-�	�	���8i���x%@��1΀�ž�
�S�e�v�G�4Bz��v2���X�.x9Q��uy�o�-W���!O��D|�zY�,���JeNG�b������]�~�V\��du���1�F&��k��VE҆��!�g����>yyN�k��VG0_�����;QR���*���W�X����H"�y���z�*�3�p`����;r&��x̂?Sm��R�4Wg�'Z�r�2�fpe��7��fA]]Y��-�G�[=W�U�}(�PƂn�$����9���%z��l��=PF���:P����("�6�x�nU�䀒���h���U|�`A���]�y��XRW��t���u� d�Z!�3�ִR����o�
7QX��Vc&.^��� m�6f�F�+�r��{l�v��ÂQ1y&�Q��eg��B�C>��Š�G!��v�ߌ��0�4�Z4�;@�۲j�)�-H��v���<��U��������׊@
���K���g�����δȨ��:��y01�\䲔�JL���*/Ճƾh�L�@J(R��-X_�Hl���Ufv�˼+��Ǯf�=g�� tt]���MdX��
b�Hᖍ��Zs���*��c�i�i��M���P�r�JC�b�m�pzL�n�mZ����S�c-϶ɬm��TЌy(�(fT��Z���yn��0l�����I5\������],a������Fx/:��M�#���z���H�?(�	��B,x�����x1�V��W��e�~�
���}�����)%�����-��ާ�lV�:s�ҧ"ut��#o�����A,�@�o[_����.��8ev�r�=k�$o�+۵�A��@���J.
�����Я������l�f-����*<D=�`�m�x���$�x����@��������
)�f�w�o	��.���D]��BYX�^P�utInj��(e�'���a��\���tu��A�OA�{��Y:�$F�C���J���H�+Nyyp�M4aKF���������� �9�l�@o�b��	�H���� 5X�4&Ŭ�?�W�@��b胺�
5	1R���WԪ*p7bU+x+��:
��Gb��m�Y�X��BN�@4l�ջ��(��� '4��@�
����=��#�]��a��S,��9,K%��K��h
-4�=�����V8�G��g.Y�o�jTzTZ���N��f�����g�wY��}f��֮GlsG>:��͆��MX���;�Z`��a�vÃ�*If@#7�_%rk�0�Tw qG�NĶ�sKi���?Q�c�yH5� 
�9e��dCDI��z�[,��=�y��%j|��|r����6�eT0n��aS������*�A4�����g~is�� ��8E8��B-�J^yZRe8a�&'���Y)���-������t�-?,
}I�̈́g�yЦR1j�p�OX|<I`\g@��hu�._�G�́�5�pC�n
�*&�<�Tmv�򕙊�;v���<�'���3���F,�*�쎷��	�%0�-|$9�k�Q�)���ۭ����<�K�w�?cUH�a�!�Pj�i&�';`�V�~��7�����U�q�/���1Ġ�H	�=o�/��%���PFF@�0���_U�֧�u�e!k_���Jߺ׍���A�T�1{L�E+I�92�7���y/�Kn�doE��#f�B�C�)���h{&T��\�!b����=_r�}qP3g�� ����g]���p6�߹�5���q4C}!����o���S������S�N����*�持O�����/"���2�2��#˘`d_r2�3p��+�=�%��M����0�Ѝ�t�j1Оy=���(֛mr�T*.$�3���TDudY�k�W@�͒�"� ���~.�$d���Yh��J��.q\߈2e����q�o(���._t:A��f4P�O�*0�`	X���f�\��j���E��Q�
k�$���M�����28��;^1W�<��`�y=�X�����o�קj�8���q��'�Pr��*u[2�;%|f�:�C� Q.u����0Q�����Ո��Z���W������(+.̏��1�:P���|�(j�]����4nB��L��7��-�Ȝ$?i�%>p���F!E�Ь$v<��9<�0�����P�����9����}�q�Uw��S�[��R��`{_Z.�U♚A��lo�{��H/��ߣӬ3���"����!Q��Aп�I��l�Yp=�^X��-��ų�����V�4Ѧ��������rM�; ��������O��]9�-M���F���1���̩�_�J}fL���q���0eQGz���"^}����C:��G��Χ�2�4���y�|��5��->t��RMĚ�ƛ��&�ȶ���M��oih�������ʦ��������.�{�x
�rWX���]� ���>��������dl�6n�+���̋!�8���9Fc��?o�1+�Q5�%��o�9�YJ�~'  K��o� ,�Qi������V��Ɛ�B����-LoSns�0C���S��܊�~���3�1'����&��vJBl��%9�����to�X��-�EA�r����@�_ca+)J�ݍ��e�A�
LQ�Z
�Q��5�d�GK󸎨�X��M�wa��R��S�g�wnh�b(�PF�sP_��_yh�A��s#/)�p��5b�	�3���a1V����E��h^5��K7�$Mr���C]䱮��pi�[��Ã���c9�z����PҠyO��W�����q5���F
����À�jm˽�ٮ���]��S5�͇�85��/u!�/z�#/�Y;c��w��E��@7ˌܯ1!2U�t����tH)/3(��NBҢGV^�&�l��j��Zdf]��� �2����G'��]�%�N �p��\w��+�q)�~��*2��q�0ۂ�
�4~2p�7=��
����3(5��=
!������R����8r�tm�҃���r�v�� �PЀ���`���W$���A�U=��.���f2�_�LI����Y��C�&����ew�m9��F���唱f����S.��� ?:�7�ڗ�^ڇW���A�,�*I��/)�6��6+���s���G~�.���c�gw��؈��^=~ϲ�m�l�k�=�STIZ^;a��j,�fPc���;S��V�/��Q'�"�&4���	]\��ذ��[��/�]}�C�����MuOo�o�ik}`�������ѫ�{M`��yu�XЗ����w�b?��T}?�DZ"	.U�ʥb�@�g��7��šZ�הU7Y-k|ۚ�>�R9{j_�6�L����+��u��+6�m��}0R�p�L�hMz�<�e��Dt���^l�=�yr� �4뾡e���Y�,�ޮ�$%ޱE8��޷^��6�t���	����h�p�%�d���s��/}��Ձp��r�S�
��0��+��6\�j�����Rϑ�
צ��>��wv�JM��|f}S�S��3M	}�|�P�JOsGց����u��1Op]����6��SM��5J�u�(Ӳxh�d]g����Q/�ϴ�@L��4i���&��
s[р�ţ�$a��A��&��Ɂv��8���M���UxBS�i9}��0�Ċyrg���ζ��C�����1����p�����y�����/k�m&e,dl��;&:v� �֕����zXɞE��OB��;�À�l�]�'�\��l����f�|�"�g4U8.�ǖ@�/��� ��J*|��a5�Ȗ��bT�^U|B	UϽ�`�]�!�ǉ� ��%떕ڌ&���
�׭~I�0�_*h�����(x�kl�_�� �J��i�����D����vC?+�!���|�����o���������3��)����U��(�V�[G�.�M��f��bn�e����QNg&V �Z�EmJ�P���4���.���l��^#��=���;f��沟q���u����D�Z��*����'ܵ�P����Ln����4���NK��8�ýù+�녠EA�yZ��X����{��:�c��G%<��*��w3�.G���%ִE�<�?����T_�^��lmi�vT�/66��?c���v�1���<��S��@�f����1�� ��&{Ȣ���r�øa���#�m��[-�ݙ��ELͶ�BA����&��;�;F�BD�_�=���1��i5&���Ā�)S������,���PD�Qq�Ǧb!�.��˯tJ
�㎤��iFi9�amH�=�$�=�V�ua9�a1=CѱA[CO05Nl(�x�P���G�c��t�i�gG�����T��`s�R�S"�aL]�7����Es���i�ϧP�T�d�CA>�"�-`V\����i�����`�^&��aX��W���J�Am�g4$�E��z�,���<^�`��B,Xg�ى����6��S͎"|v��ܗx�n*D����4$�f.Q�_���j�ԚԟoZE�\nb'�[�ٕ�M���(��3�0,xM-c챋��yIN-.O��M ���Ua����?�p��|V64�6��=긝�0���:�v�aw�v�:��,	5&1����@#���oNSah�B ����=1w����So��
�5Z���q��1�5�� �&v9����Mi5�{��Ȳ�P�5Յ �"�4��y�hc�%�G���< a��W���Z�h��>��v�p�M�]�d�Ulf��c�����@U�Ab˵�J��&UU�P�sBV�+��6�4�-����U�R�_zE}d"���S\8_f�(-��V�\��=�� _������t��|���#`�
UNBdP9��^��W�ї��ߐ+=�ďYO?-��!��c�X����W�9�Rw�D[���0���m�e:��̱ld�ږ�j&BîmCse����9q^�Ɏ�у*ߍ��+{_�s�<��as���y�#Z�����)۰�i�]���uS���&�Xc	�Xε�@�-\��+_��)
���<F/#VY�W�*��D	����}�n͎����q>��Gq)�"L�H/^�MY� wM�X��N�h�D�,�%�����oi�R^U��V4?�!B���L���P`�D��킅>���ס�$�B��2��ݝ���>�lx��h�9|�)�� ��䉛���N��
^�ǜѭ���o�+�;0l�-D�r,	v����X	Hͫ|��uSDht卛cʙ�F8��٦Ң���@:灴��Jf��?�v�{�Yv㶎z���E������7U���h�P�&;]�'L2���4[tV�&��Ľ�<P������P�vӇO v,k|��57�l�e֖��Q���֞ښ�]���T��E����2��+-g�����
�c鈕��w��ε�ǵZ��`��*����⟊�\��@��[��Xk�C-���L��`W�a� 	Ğ���E;�)�3~l�O��s�y��]�����g0�R�\�yw�?sV%&�؆����2�[$󇲍_ #����:��CBt
]�*9������'�GC���'`:��J,�3l��GR�����tWI������jT�5g᠘�r�U-��E�X{��*+�2@�mh��Ȕb&?zJ�O 0�Z��k����τ���L��[��Pv�ۦ�6y�3�1����|	�d �n��i������k����!`�Q4�푒8�O����sX��	��xl?�����@fV��|�|t.�r�j�@$��/"�h��ؗ����n^S��%�ϊ��|D��u��Nec]�l,�	�WK�N�+�E����ޅ�nb�K����5�wF[�c*j���a�!�u"t2��t��������}$S��0�?l_�v�&���\����^?ȱ@�&���0���hA�GG�C]��)a��������FJgh���s�A����?�F� �x�C$j�${mY��&�<�UV�����Cq�^���o��c�5ٹq��v�2鯇��F>qqތQ� V��9V g5GU�rF���q��o�D�l�V�����|�Њ"����N=�� r�'B�$l�j)�P�o7�gi7"�ׄ����i=�1��4� vߟ�,.I���u�e�N��JC~5�[�ߙ��WB}�۵	B�	A���fh=����怮��1����F�V�hR�%CN����+(�z��G��`�:/������$+25.t_%x>���w[���IY[m��+��UY�Ēe����W�&�����v�.5�LaنE�Y�5��o�X� �?A*1��Y"�i�P�E�q�\��6����R�h��{���M�rdF���<�ǰnt�O�f�Ay�|����s�Zta0���>�G�;�Î{w�/,�����J�ׅU>E���{#�06�ڗF�ĵK�O�<��dMqk���4��
vAQ���IC����9����܏��\��Os����+,@sxZ����
]g��&��E9b˷W�~�(>���_����hE��O%$-y��2qR�C��z%�87����(N$|�J�z*)�o�� hi� Z�U�ٸ�[K���J_���dn����W�m���!����$^�B2��7�gL���@�nF�������I��s��;~�bۈ�>\�'O��!ĕ����2'?w�)2语>90�I)b�E.#�_z:%8l,���/~T$���PxS@�}rP՘~%�����X$1�e�P� �Y�$͗���=�P̧�K�|p�u�s;�)�26�t�hPg�A��On�U>�����w޴�T�YfY��)/�?��Vt�n]��<Z�@�����6ϢV���K�C����Q�JP��k�11�e	^i���Ŗ>_��*}nG��{p�%>~�ٹ�iz�v�I�?P�s��O���̸��sh}9�U�T�K/6��� ��htw{\��W����1a��e���LJ���zN��\9����cO�)�X\ų@�{\G�:�ڪW�%�JTǰ��C?��=�����[��~�MU���%mp,u�.��٢R(ˣ��[ȝd.G
L��+P�Y]�[�������Lr�r�����*�+p1���nV3��?*�R�zK�p+��m��}@���MR3]����$��c��F7؀�?�edz��R�e������;��������QP�1�.y(��'>��ưN��}5[^IǓ�H(��^6�ĽH�0ܣ������1�x��."�L��>zZ&��j�����\P�IG�)�cVX����d�K��������oҪ��SE��t�LJ�(K_��$�{D�1!˄����t�yԞۆ��{,��np�����p�QXѧ�h��{��m�\�w�e��k�V Q�:�sl��VڥS����3���C�/�姛-XY3���ۚ_p���Ef�ls#���+a��Xe�6���U<��ج<p?��)�FJ3���</�|�����Z.��ҕ?aS8mݚ�24dΫ���=�2/���u"F��� e���C{�"d8#J,�k��M����^Jz�|ξ�n3�H	����^^�EÚ{!����f���jO`��ԟ�$C�۠lN�����:��y���X6� "���>U��c�Zǹ�WP��0�-�6��^P]۵4�1 b�RhR��-pi0��WU�+�ź�f��=�U���z�oSL��-��� ۛ9v���ȼ<�򙗸�:��q"l�oB�ٱw|{Ykg�7�$��"�n��Z�[��]'LϹna��&��7�⷏�w�ߛ���)�A���tN1}�{�v���'�U�^�W�̓ء�8e7�E
;>����H�u/��Yl�W'`y���O�6����W��6��i��u����_���>T>��0&�������kZ��!�XCNA:
e�^mb(�Z�9;���}?F��w�A���{7��~(П��Q	������e��͍u�[�]�$ s"]�:�kBf���i�Y�����1=r/��x�Y������au���^p�a��/e�{��7B���&S�G�S�dI�*�����o�Z�I�'�i�Ϊ�	[���O��o'��ύ��N`;�SK�g2�jM��751�!K��\Y)�j��� ��#����tx/���l�\�O��v����DB<
�v��	\H�p��ո�;-k��P�Ԏc���T��NF�T��4�@�����pH��/Ė8y�������2.G�6���G�~K��ͧw��	�Z# �d�Rksǔ")�t�P)�##�� ���?�ꂠ_����J��|_����:���t��AX��P񤓋j{����~�Ս����(YzwOѧޖ�Glq����k%�Ѯ7��-G���8P��r{�Jj�$�mk叨z�?�w�|4i0���,C7Bƀ����WE�mӛi#J���ʋUR|�I>#�9,˷�;::p�e��Rj�;��;�u�DЀ����>O��Kr��K��^I�^���<&0��J���q\�b�8�MM�	�5)��\n�ǲ1JFuz?�`�'��� s�-���<�7�_4>�O#��{��6-&���sr����>j�%TY�����v�L�]����D��㳢�q����/�E��ͦ����Q2����d��+m�S�X��;�ؿB0E�a���um�w^u�7Þ*y�p ��\��(%��0X�'GH�� ��'֤���wa��Ʌ��C�����>µF����S2��44O	tǟ�7l�cL�1uϳ{C߸��QP+*m�Qq
I�3u%g�Sy�R�{��o�?f��KK����2-� �]E5츯S�,���i��)�T�j�t(3�����̟�C���.�ب�ˇ(]��!|��e/r���e�~��y-���/�_��sOn�A4��Y=�ҟy���)mv�%~/Ҏ��p�Ez�����Z�[w�����i�VӍ$n��	\Z}0�p�������G33j��Hh�6�����8�no���H��R�3�&��+�!�(�S�\"T[1oS�W#j� Z���|8�cɝv������xx^�^�NX��tcI��.�@�=Vjb�O��:c�U��W��Mq��C��1E���������tX����~˙��Y�V&���Wܫ6V�}R�v7N���@ ժ�I3�"#��!��:��k�2	P�*����'�i�̓�}˶:����2;�y���1ݨ?�٧ĪK�8�=�$����,�%;�X����g�xS7"��*h��Z��%�T��!�?��8���j��;}�Ȣ7v��@��:F5���S�62䢎f�q��|�Q>��|�Z�9���vO���
}m&Wl���{\LT #?|f��i�vt_�&6U'�؁��~G ���0Gg�?AK�%��{��J6��c��ݣI1s�A@�ҷ����|�XP%���b�K�R �����Y�c���z���	Z?�z�eߗ�kz0�����NL[������2I���v��J�O�7��sU�������;���4�D�E��
���}�(ZZ�E#��7���=�����gſS�P�%��L�MČ��X��E� ���>��Ȼ7\ߵ�t�_�Xj��Td >]�$�-�˼�ٵJ�n[}��E!�*s��*���\2a_��|R,aRz_�;o�m	4Z���$�J�b�>0��o�(u_h;D�w� ���b.���:f�'�O�Q�e�����<U��ZG��~~�ޝ�'�˚x����.ٲ�pq��y�à�Ƿ����F�.o�"~�7�L��-<Ѷ�����t	����ֲd���_��?z���dl0��X�'J������<|���	�����6Zn8>�%�f�F�d8�x
��:�v�)w9
�ۯ�w�
M�µ+#�,��	�D�dܚ~ ]f;�nJ�)0 ��.�TE�+�Y �tE��:"��ɫ�gt֪,�;��6� �(��>����{c  Qs>G	E�M�!��kDg�ڦ
r��u���'�/ψ)/���.O�q�Jފ�4��ϝ4"���^"w��.q�o��OˏUu��s�@���J��[�X*�Sx�ʘ B%�����3y���lq��y@��^�
��8^j���!�����*g�l"p�4�]G/Eb(�%l#w��Т2�N�n ���1�p��?�q��Ӝ�@�U��8'f�@�]9��O)�T�9�:p�?'JE�3~�>x_#�ɌO�@�~@hq����"U�z4/�-��bzGL��V�0���� �ݵݭ�Md֔a��i����C͓8;�G|� �P|��p��S�F��������B�/NVŎ��b�Å�"�?6��rMg�y�Q�� �֟��M���Dnf�ۇ����k��B^���}8 �Y���:(���>701t{��J�4�-`�<0������Qڀ��=�IQ�-[�cm�3�����ICM���\|�-r#D��1��݌ U0UYCXdS��)���6��̶�)��Ǧ����َ"5��	Kꌕ#Y�|;d�f��\�����n�SQ���v��S��#�q-�U�Wr�eJ���ܢ����x^�g�I@]!�mcpYq� �v�S$?�>H6k�~��+�l'q����-���hJ��'P��Y�ͷEV���#tF��}�ڿ���(��L��bk�ՠER�܌p�^�>���Z!븣,�jG��9�qlp���͗7�4:���U��SK X�����C�	^��Q/�B�����4���q�|�j�E��]�fs��(ë�|DH+�e������Z4�4� /��	�V��G�^�RV����d"XQ����Q}��x��:ه����<����Ͽ�{W1�8��ߐ��i��Q�O$���O��_�%K� �m��t�VI��2��Z�n@8%�������S2�υ���F�?I�q���uwKc	������M��jh�N�`��F8k�����h��������rJ����X�M�e��OЈÔmY	_�o�,�׳bv�Ÿ����-�g1д	_s�i��ͪ��9�1���`p}"D��z�/I�C�����FRCW��D�tٓ��Pg~�$�C� K5��N>��ưM���Y��&�'V <�ڗ���+�A��׮N��j9_��6>�W�9�3Q|�>���D:�����B�X��Q��i�������rg�z��v�i�>�Ŗ(6����	^�瑝�:�9��ك�/x�5�hM��y}��0�qS_��w�=��ű{sr��H��91�w��J����y��z�dI��F<���X����fG���7����l��=Fk����O��C��ޯ��G^u�HՇ�7tvUbW�N��K	�joD�b�yLQ�sOP�D�ʱgbvL��~��	�UV�N!�[X=�8� ¥�g6-Q�F���������V� �Bú4,��੿%%�mV!����{�]d�oQ�è���(�Ty��{@��>�~S@��nB.�KYg�ڮ\�w���Q�(�3�s��d9C�ck���dp!���ފT��L&X���%��O@��x/�l_;0���Ώ^m�@�Ȗ����7�XW���x2�z��d�.����D3���N#��Ô�~eQ�t�Bx�"0����y�6 ��`�q�N2a�
,u��#�q%S�n͹G��lT"����T�S�L���3��~r�HC��k�;���s���Z�=�`=kWz��n��?�q�}��c��9�>#ڈB�]M�}u�Z.�Z1c^���k�T�J�H0�9TkJ�GD���7��U���Ȧ�7cʪE	�z����nՒ�$5��m����9t���O̵�dh����A.�Q��'K+����3��Us�}
��X��ӗ�0�ŭ�I�R{�KC�����$趄�k���Q��� w��@F�� tF���?���X"��4� :'M�P�]���������B_Ʀ�.���G�B��j�=��&���{֒�s�r˨u鄁�OҺ�m&J��*vR�`zo�����(��-ZN���c�b�ۯ��3L-)�������jʗ}��A_r{��E�GK��r��S�Ѣ)��> 6�}��#E����	+�17j9׏��1AFA�
-!��U$ɹb!/"
���Yn�rӎ
c����gq'�d=�I-�W峵�jJx��9?T��i��8�Qq��)�Ǧa���g�� �'���7�ի�N�yN�w� �QJ"E����j�ӣ�y�v�ˈI��N��U�((ׯ�ѵ��@�;����TnD�����ng�D�uH#i=I�ȣ�Տ�K���E��N���A\O�� ��{K�o�`�X��˶o<�6��x�0�@��8���L"�n�K�����K���,�[��a䅼�/�"�ՑB�Au���I�3+wh ������{��j�c49�!$��c�U<1��ِ��_�f]���%�<�1Q� �LNY�K-���:����pu5TT_)Ƚ
���ʎ�! 6aŇ�7�1'r��~�>�R�K����-���G��m������M��@���K8��츤0�a��?Le	u�]`���
�<��\�7���+Zӷ3�L�����#�a�"��߅���3��?E��ׄ��i5������ڬ�چ0����Vn���n|ź8�_Y�G�P�n!7|����&�kCڧ��Whi�]ᦱ}`텃߉��ǹq���PR�[X�	]�5�	�K��+���
�������﹭��z�}j<�F0�:1I��%G�-:���� M�nF�\M�d��$�;�xK�� ��4�֙�=+h��,k � S�ҕD� �.�s:����e���ۄ��S3[$���O��l�`JSÍ��>���n�jć;�2|�d�5P�wp^�p�aǧ��~�L�`Q-?Sϟ�����@i	;~���nM<���TW�m)̺G���aq��NJ�@�(u%�fU����5F�xNA�e�W�Ǥ�y?UN�8��J�=����p���{�d����^�t���TI�P�G4�J�:7����X[������5� �pd0'��V%s�G�4.{\u9�S����N���iw��<V������ݞ�6��3b��z��Mr風Mŕ�g�5�Q9]0+�8�vA�U��������&$-'	>ae;�?�
�桑锷|�3�Y���=��`�M��4�Gzܜ�l�����M���R��-ҧð鈆��<Eۖ����kӚ)8�՗������X��w��6g�(fP5E���U^T+��/�pve�6��Vv��䧊���\�8g�JO@W�#��DF׍��)��uO��ԋ��Qa�9�j�x��<�L��>�|���0��/==ͼ����,�gLurx����{�	�}Dƈ̯k�"S���gA��呈z\$�����������04*����D�s�����ϸ��Eお$J�M>s(�Aގ��]k}Y=?dW�@D�a�?ZM�
��H�%���v������inh9�?8S�o�c�
���v��:�.�Y�E��d��>1W��-A?t�:!&���*�5М�[�81TĒ�O4O*�R ~b�����jc�|{�223&K�V+K�"Ӵx�g���4J�|�����T��T�.9���u���g^`�\ �� �� �j�"ݔ<�]��.�hLw4�a̳��(I�����>���`��<�Z�j��	]P?��K�^f0�A�'#8T&z���	V��+�.^���	';��i�M���g�ºwͺ��3},N�����c�-&���n���4Go��Ӗ������iU�mW�@�9/���[l-��:5�cb��x���)P`p�@�������W;���r�)��,|��� 1�%Fu�z�(���'�xhJ�/�bG�
]n�$>�f��H�:����<y �:�~�j� �)u������Yr�+M���bU��h�o�X�z+��]���Q̀�L9+uQ���Ns}�L"�Jc��aK�n�%=�YV�.��$_�:�q�~���<;4�n[���8Ap��vz��A���d�������n�W�3]�DX�
48�5ͷ�T
��`���Gm�p�B�;�x0���o 7�Z"h�'��B~q�a��Ħ�����"(U�Q}�,U-s���dB-<��4-{'B����("B��4"l�K7C�܈����f-��G@��X}]�\vl���t#����!�S�³�e��:���zM����eZ]��am�č��������)�x�^c�+`�D2w�F���{�N�*'�g`�����"֬u�M[w@Z�~�`6�YNФ�" m����`���e�Y�������z���0���s���Nk�f0��}Eal���	*���=�8�$ ����j����F�Md./��>��1�$ �C��( ;���)r�!+�v�Kۃ��ٲ8���bn닷 ��}')�e���+��j4�`oI��)+s#�>�(i2�;�;4]y!�u<Ɩ�jqd*�,>���h���t�J+bs4���_�$�:o��l$u,�6�Ɯ�_�ۮҹF�T!,&����] vX����0�b3��0V��h�r>ȸ�рf8	"$�{D�+v^T �6������-O������V�����E��2�D�x����3d 3�zkb}HIk�����p�ƣ��ųi�(n�y=<��"+��ٓ�P�ͦ��I����������؉��q~Dp��9_��Q#�:��Yb%/���2����D5>��-]r��	'a� ��2�*��a�Jej#H��/Z�V]�ܒS�m���Ƚ���Qd�^�f��(�B'&@z<Q�Ŭ�e}�3	�OQ'{)L�焫=Ѫ�b��
�*��K�i���%qGy��w�"V�!�R��bp��8�@[9�VzWO��h�g<)jD�i����9�U��0�sE�O��R��p���'E�k�]Y���8J������ !U���!�2Q�w���'����,�W�r2�3��w��P\nB�>�����7b5�d�B����Hj��+R �l�ہ[�dKZV�/T���ޒCz:����1}��mݘ�9:�V�+~��7�6x+�!	�&�;S��L#�W�l!���e�Ў����D!'ԄO�x���s㏍�C�b�`$�V�91-�^�|����ꢫh�C�� �����ntf�d����t	�8��e'���F�[�׮��ն�S�X	��L�;��8���J#3��-p�ϘW~LFmš�I����_��x��zEE���%/D�:|g����!�I�lI�%��᧣q�5I��$V~"*v�J��ܓb���&z��I�s]G��0@�- ҥ��`�$�.j� �<�֗�*���Jh�Uմ���aԛ[c�)�O>��j�8����ᄔ�?�)��Y���'xg����1R��Y�� Q{�8Πf����-��� <㴲�)�dip�l���'y4��	3����N�:Q��i�G�;iZ��7��@�k���-@���~������;XU�S�V���/�i2��j����٦:��b��4�<�n����!~5k
o��N�'��.�'�d�\٪I�i=�x���mj���X�qP�u�	���f{A�d��E���dm��{�{��|>�К�U�hmD���5�3���%�{6��	:�~B�օ�x����oQj|:y� 2Z�+�T����ʳ�-�d������j�$r��L�?���|[�wvEc�x���$P�1�cV�YXl_w���%�����;��G�!S^�z	/�Bl����?�W�0�n[��	ɭ ay
���Z
h�\��V9ԣ�{7
�ن����AX��Z3��]J@	靛��;#�;�7�`�a��E�z�Gac�,ڒ�ؔdf,�:��i�O��}{�Nkb��:�|���ᚹ�b�v�]�n��������F���-�[]�ڨ�ΰ�@��gE�b(��Q�ƽK�^�{����Gc2��wT4�Xf�b��NU�[���	"�ވ 8������
#KCB]�O�J=+�"�3��ݨ��rWLge�3u��Ek�N� ���A��ᯄ�Ղ�iĔ#�ρZ��O �쵓-X��)]���C�	V�S��i'yb��Tl=�GݘsC�o��6m
5��ٸ�w7�hZ�����=�V�X�_ͥ�'�Xk�����ʫ�=�v�&hmj3;k�����=D�w';:y��Z������4e�����Ib�/�.;���$������3>�@�r�x��/�m�j��pJ�e��_��%:���HW��5��ٟ!W���,�ƈO��w ��7{K dq�N�$T�p�q�&K��c�s��f�$K���0���=�����U �Vx9�y�_�
v�Dg=g�S�?G�Cn���}�4�ON�D�P�n��y�=�z�ɯJ��RT��y(k����u���`����{H��ڗ����聓J��� )���G��Ό�#��ֈ��r2Mho%Ӗ9 ��^tfv�}�<K#�ݓ��.�D��U.�\Y��X���_��:]Z��b#;���VLi����y�n��p?O��:��k�g.�0N��2��I-���E֟XϘ�X��dB`c_I�+��$�T��\l��H�W�����y�v�v{R�Q�q�)��=��h�@��S�<"����:�3״m�^S���T+y�9��E�.����������d7�b���N�v��~ v��?��C�����oԥ�w�b҃w�ƚ�[^D�r#冓���,(�6!bĕ_>���~���J�-���ȵ�\�m>�d����M�d��%��V����3\рD�S9����|�-�A?V��� �/�ЦH����K�CH��K����֣��~�x��4d)w�!�Y+����i�:p`N�|���U_7����lzY;A3�Q�3�{K��Wi"�AO�ui�8�Xd룽ض�%t���Đ?V3K�<Q��25�����1��~��ag#�R��OC�s7�ģ�$8��%c�d]���$����:
>К��U�����TȂ���ۚ��X� �z#�U��2	�9�N�:,%��)F����M�T�͎
b{�|���[W�_J�7=tm�i���C�0������v��cC����6B��|]�� U��s҉|+��s>��'Mk���\�I!��q�L�}����p�v��vY��z�Sw)F�#URnA�#�Е#9�.^�(�W���}�|���$x��Ii���B3\-[t�?��K�{�tL���o�/����pl����D;]��z�������l�Az)f�Vl���j! �gh�0��(u//����6b�q�h�\t���i"���B�LҴ�h����Y��mԔ�Z�G��˪����]`_��$
o����(m�Y������
���H׀��CY:��ᵊo���/�K�r�Ñ��Z��Q?����R@�-�dg��F�����^���ts��=a�۶�8hV����=�,�t?�M�"A����P��`cx=�oA���dx��U����hg*����\� ��,qYmO�ƝO�B��K�,��Z��!lL^����ץ덛n/B��Y�dG�>5];g�Յ�l��>O�?���mxlo�N=��p�6k�U	CTH���$H*w/4Iq��/ě2SN�w,��מ��F�O��.��*6��̇����1��{'@2�b-{]��F�U�Х�ox9R��-<e�{w�s�����_q^���k9�w�{{ɪ����%C�$:-,[Q�/I�X�IlB����]�O���o4��	���-�r1�xG}}����;ba2��-�=�2���n$�����ȑmD�h�Z�a._q��h�X�������9�vr�怿��aMS\nA��ܵ�XNjK�U��uY��*̇�X��;K��H�G���k���1UǊ�|�F��`G_Hk�(K�ڶ#��E��gY�N�nt�hK�7���Z�[|��3�$�X/�j_�V\�w�J)��`�A߫�Π�z��MUY+�8�Hy��?5��;�@�(t��Ez��e�@F�PƙB�����"qEU�@4k�z��O�iLD�5�\k��$ʯA�l��S����?����f�#H�B�Mܳ��V~�ꭲ�b5�w5����A-\0c0�<�d0�#�u؀(7���)4U��N�^�՟�΃��
�Q��'N�T����>��Nۦ:AMêg`+�z���K&�[U�\彯t��j����dLқ���Q��;���<6���FF�Ġ�ϷL�2��^И�ɃA(��,��I�RU� �B�Ĳ+��VRɣׯs�I�ppԨ��m�d8N6e&~�mlh�y9O;��N0�m�>��L�,*���½���g��7	]�ژ��h�Pl���c6~Y��蠂�@�6i��mi��$��W�E��~�>�&nk���JXr!���*&A/ј�
�p%��
�,d:BJ�W�
|<_�No����O�{�U�㍔!]���;�Y;�O�D��z�4�'�c�i`�Z'���N֣��Q�Wc��]�@��p������bVc��T��H��&'R1�'W�-�#�]���R5{��t�vE�{�����˼�y�0��te��y�.����4E���Au��˩@���� �Z��)���U�@!0=�'��0d��Ս~�/y	�q�F{���D����E?	�뜈�*�7�4�� ��c�{�2 �$)����q�5&:��b���V;w����J1�2�Z��qG��S\X��4�@������1�J�����Z�9�*�ŝ����K��t�v��f?�/{#o[��(X�T�έ$��,nh�V�l�� ��bF�gb1�zo�=�_1)z��r��Y�[�d\@�C��ay�xY;�>匱�KA8ǒ`���Ө������{�޾U�R�v�+v���m�6(h�$y�V�y'.��ܑ0���P������(yǊ)U:��W���� #��7�̱�V
����~$�\G���e����veM�B�Iw�%�S" 2�b
=�n���Lu.��e�8�o/�3`2bH��S7op*�j��]�÷�c�gִ��i��f`�-C��)��$�Zā7D��%�}mP�V�\Zh+;*P������0J���X.�.�Yk�����GPK��zӦ_a��˘(I@�?x��-�e��u�ڴ�R���8ʧ�<�Ķ"�g�jB�u�<+�`��L�k�~g���?{�W��m�5I_ر6c$�U�Ʒ�7���X ����b�"u	Ɏ�k���bj���^D4Zw�Pj�i����jo7k�O�Ll.�ݛ�B3�R,��s;Ǽ�j�4�w+`���vV<0��E����*î�;��'�(Uas�3@6+��P,�r_�������G	���\��n�� iz�M?�,�M>�bY���r�z/�rRܠ6��\3��C(��9���z�F��@U��0F�`�p���Fh���[{B��� �l���4ד�Ь}'؀aX��2��Q�8�_�:��.��e�D\����}��@��ȎZ7vBu�p��Z�ܳ�wukm��?���nL[��1f��(ik������˪򿕤S��ɘ!�*K�u6�25�^�*d����m���?bYR�Zt-�R �?�-��s�B
zr������.hzd�ԆU�8`d���a���)&ӗ{�LL�C�$%�#C���[jɅ<?�6�D��M6�.(g�#Y'���>L ����:�x�;�!:��c���H{�I�-�y~v;2��,��eW.c��n��C*�ta-/�ck�X�ύ�����À�<:~���Р��x��qqRo)����
�]�. ��sZ�>i�Փ�ݼ�M P�.Э2�h�])~�o,�(��w�,��J�M���d#��F��t��7d)"c���q( [��;��A;<C�M�� ���)�t�����Pw��؎pJ}��J�w��'p��!Vuh{�X����|�>�I���P��c�.��oZ��:��@es�C��;딿1����m)W���G�r恱
Y7�Use�w�X��Cq���X��T�7j���GIMѺ,�B�c3�K�Y�^���(�m��$���<yT�P��ƪ1�@�Y Ir$n$��
J�-��~�J�>��Sh��r�/Z�2�O}�=��Zq�DUfI+i�9E�Γ����cb��;���&�{�d㚂����?4�:n��zi�3	�}�ff�?01hTo�U��6&Q-G��7�k�ReD��ؑ�g�P"\�<�6�7�֗:�yJZ>�*�V��LC��9,��J/�w�E�����x=$��E�H�d�F�f�!��A���(���c��?��&-�>n����#J�O>V*�-�o�r�겸 �@�=�R:"6���C,
�.l���mH�3�1���W(��'#��%2�8u��R3� �b�?�a,���Ì��d��o�Z_�_�����U��!;�O�ˊ��kl�cԡ!�v�q*C��i��F]'ra�3fo�D�D͝I6g�=1y�	�}ܕ�7Ԣg�8��Y�tɊ+��S?F9��)S�M��'�r�*L��X��(B��	w$`�U���q|+��~� J�ݙ[���]�2�[���g'>�m�Ga�7b�i�v����k;�����0�@(�[lvS�ǚ�=������
'�P��;OC?��i �t�+��O�/�}}R�
x�tב��U���j��i�,1�R�i�����E3[�������x��3�޲��6�_n�OO� ������#s��9]����r<a#�k�u��O_\���b�vI�!���� ٨�u�p�z�8כ[d-x�a�i�>" �&M�/�Z+�0N@nf��9�\aF�7e���բ�v�#�B-���*�ϣ�@ѧbX3�J���O�4�9���crb�gbۗrx	< Qc��b�t��@=�j/k8=d���g?�StN���\'��H�fv<���ZEO�d��}���s�|M'���g�%��� ��ѣ�����hB�KMF��N-d4�2`�Cл��{ ၬ�9�?vß��y�a�Ib �Pj[x.dkB��ĶeL(0+�Kq�G��d��zI��w�}���`LL|kKL%FW@�0�V�^L@���*����G_\cU?���g= \k�q����N�5T��F2����i ���R�"7!p�ƅ
�0�B�56	)�+��!	{����t��{�0���[�a�R�Z�n���= ����.g���d� 1§ �'�P_V����'�ң�l��B�p25Q`������S͗1�r)u��.���Y��Jc�K����"��b�ʒ:�d��G�sMS���|�
&f9����[@hjR��w�]�/T�ד��B_h[��	�vJ_��@��w޲IV7��� �|6�\fb���{m�q���T$��?���z��aV�枅��@��Ƣ�w�+��ӄ�U	�D�˦�?I�2���0��;d \�d0'��9GD�0�����lW(lv(q�ݾ�Ћ%Kc��tRF~�Ҝ����i@��&���/L[/�E�|=^RSn������ �Իۚ��g�|^�l1�̣���U�)���ж��1�����B|_��">:��F��} �W�\�n�v�0�|8\��m��ޝ�Ӷ9�Ѯmv��T_n��)H�v|��ޟ苺�I4��Y����.=�+��h;u��b�HBx�s� fk ��;�Ȁ��&��/ L󕚵��F�!Wcae��X[�{�CkI�I��,g�" ��x�*�̞?��kĖ\��Uq�k�>�VCSvp��M���6��~����o����f~V�F��K�i����r�[^CiZe�5m�?��Q�ԣ
���,�S5�ů�!L=��X.CH�X�dL@ K?�r}c���59�v�n�3��Qkyi��w�������q1��������<�C�wk��f�ua�J��e�����$��!J����n���3͍���-�8��Z?߲��#J�G�Y���e�kK{'J.����*Ϟ�5���3բ	v���e:��^�;
�Hhk���4��\"�C�x53���Y�ϑ����؟%*��dןs��o;E�R��D`p��K��C����IU�;e6vB�I�tP����^�(1�q�d\��آSJ m
���|ɀ�; C�a�v��E/���sO�Rl^���UJ�u� �����]PTh�<0���wa���C���,�wA�ayqj�����8�fe�c'�@f(�����e�ߦ	�YbTP�6�s�:���bgG�^���9�4��v1./���VY�a��Jͳ4"�V޽L�~Չ6PnJ�
8�Qï���qA��v����
�F�p�eR.����(����NA��R����c���	r��$����LCs4�u�W5v��s�jG�v�]L*Ϙ�����\��R%zS��jjYhV� |�d�ta�_;i���p~�C��]?�i�O-����k�������y��g�[#y�n��k0����u�d�KN� �[@-�_��z����X�ۖ^?��E��f=�?�3#;��:�hWS�5�N��)wI�YH�S�acϫ�8�����I�2�k�G��ip�J<�/�|q���o��@�I�
�o�R�7w��&���Q2.�-ͳx�����~��f�� *������W�Z� ��u�P�����x!tYk��~q�·�c�cM�}�}-�aI��2D9�G�������6ĵ�b�Wj�_��Ḥ�S=%eؼv�d7�y_�V^_h��B��ѹ+��}��Y�-TFNw$����ơB)FW��}{�
.�Hqw�jUr��]W6JR÷����rA�R��%�*=-,�\4�}}'��m��m���3��P�x�
��?0@IL�J���}̸c7-��'chjC
XCE��)�!�F���ќ�M�:��('ׂ���t��n���:�<N�M s��"L|Iњ��x�kl�*/T��c	O��6���0>�1���w�d��d��!�,�7UX�E�<��R|�J�~��(wu�a�b�( ���x}���)�R*ʄ�;���5��Hf*�q��!GcHG��l���֙+苺�״�l���<�����ݢc�P��"\y^��{�/�oV�Q�=���}D�a��2�Q��3ۈk�TM1�Զ��v�2���C���<�ފ;v6%;e/��X?2���}��<o�*�����?p�@W��Z�զRRi�tʅ4�0�M	����Ь�:A3�	���X �y�]>�c�7�J��؝�k]���>����ď���@�%]^��r�M2g7�>��+���[	�]���?�C�\��Vs�j�{�ֺXy��HL&<����O�j<��M�_E71dh�g${"%5�iN#��3ڍ�a��&ԝ�Boy�fk�b�b�Y\�̹xэC�4��񶜇����O�����ʼk. H݆�8)R0.��y��'cvj��Do=�?ŏ%,<��fx6�R�a�H��j���p쉄|W�9"�-���]���61v�#��^�O�qr)���nH���BS�����5҂4w�P�<�ٞ��W����}��=�|�xG��u�bh2���c,_8���Kd�f�j&���·�k#��+
rpطI\ag,�*5�6�)�+��#LxO����!�2X�J������C��!=��10|�|�k��t����K۵��4��ۋ^$QB)�]������vp$aj���S��;qK'�S���!%wv��
�A�d��e��H�A�Xt�gQB�7�c7��h�O�h���eZU=�! b��6X�aQ�)UȨLS���Z(.CVw`� �?Ш-�J �=A?���\춓hp5���:@�5j���,d� ���0��Z�|�V�B��NZY��W%
�)V5e��Խ2;L�@B�c��۾�E�70!��1���B��;�{S��:��N�:����!��C�'��O��(�y���@gY|��W�V��6BX-��{�Ok�ʅ�Q�xC�I�k�G�Q�1~�#CҖVw?D�$Fz=�9br��\:�}5�좯+��|.,T����K�gB]e��?���SO_���S�@jl�WO���{��N�<�M�?�
$�UjV�;��7��H���V��2�K�Qr�;�	]��y�4g���ܮ�$�h�_�N����R��Y��&���c�#y1��%�4��7uO�U��`.�3���%�!r � �����
�,���!�r����-��abC�Gks�e��8��,�W�L��Y�/�|ů�_����liQe?�x��\�������ddB ����#�?�>������)�n�� �+�|X(XܧM"uƽ�\S���������|H���}�E���ǘ���B��1��	K�v~&��&���w�$bw�M�S�uv�D��Z��4�~hk�6ƣ>���1�M��"[�XC!�����9��?����d�b|2�(g�Y��U���/6�-�F�f��������Ȑ���l�T�س�\r��l�#�~ZVׯ���z�Z�;P�5���g"��zWa �1�O�n��w`�NSu�s;�#��X����=�0'PQ�5��8�4�w���CŲ�*��.��+����Ɲ���Q�_���.����yx�eV�'d�ase 	 �]��\�D�b�3� 1<�x5�!���'�|m��H��d��(/w�o�f��|��V���p�Yw 0e1U��0�;��Eb��c�:�3�X�ف�Z�VQ̢6:B�e�ֿ��:KG�����d��gr�u���k	�/쏃�����S����[���'���!�����-r�i~�hTb��]'O��,�g�}�T ?x\��s���̘�~�/`�1�:����WS���T��Ǹ��(��E�<�``��P<���k#���M~T�%$c�~�.n��e,{Ϛ(�%������VvU�k�
����${�2���$�67�9�&ϣG&n�ߙ�<�*h�r<�C��֞��$Y��Lw����u�aC��ej5!�妎v|Ҧ�)D��15�2oo0~*��Jp|}ES��MQwg����m�c��M+9��YMX����(J��U�2�~��?����6O��'
C�z˶��L:�>��b���IA�XP�,ُ�����*��ty�]�og��� .Uս��Ջ��Um�ij��%,,��؛�2�I�
�o�')���O~��!�"u���#u��]�g��P���9�%���^ˍ��$�[<��w^caw}�JX_�٧�Y�{�x��tʞ���*�i��N$G��9N"yc ����J՛���N���^����|�m�A�G�?�aa3�'^����cڹ*�򍦾+s������cM�X�ʀ����YpwK<�������b"�#�Q��De'
�c�C�r��Ȏ�s�8S�<�%;�te,&��a�҃'_���<�;�n}�D]u�2-����T=!���sUR��v�S��B	����a{SwJ��J����CZ���3)	y�Խ'�m$�`����4;�
��6�Ԁͽ���$&���N��sEFy�1�GOq拵��íw�0*����T��*W!�W��V��X$�PAq�\/������A�k���둽���t�F�����Kt����M�*���U��!+	ԗXU�Yiw�����U��4��F�jd�Q%��s�ި�	�j�糍�^��~�Pa�W�Q���P����M�.2WӗsS-�DKi#��uQ��}�<�Ex�}'p�>����v��';��>B^-��u���c���J�����I��E@Bɹ�b�`ҹ|��0H	�o]�^JC��b��lR������"�t��TY�:���՜��\ֿ��������ƣ����9�LH
�6�ft7��-i.�s��Ng���W0��m�X�A�J����wn�EE�0w�fD����J�5����^����6�%
����E*�@��qscF�i��)�&�Iw�n�ᴫ���=:1F]@g�E��-�� ��>��Fp��Î���G�Z�Z�P�$Hӿ��??W�Y�>͍a��$�Q&�����Ψz+[ðϸ�H��6hw���LpW��s���&�pŭ�c��{��UV��z�w2Jν�v�V��r�YZ��V ���i���I5���9�A��{	p��v�,`d�W}�ɀ\�(�4P��H/��Gn �R��~�-��꒖��9���D3������s����{5=�0Gs~A ��q��)_��C��MX�A9�?ko�ܛ؆���?�������)�X5@w�mwV@�p�*���	�nA�CϠL��ڥ�;XP�mq���{�ޒ�c�Ù0D�Sn�o�8u@�ݓV��[]�v��Z#�1	e��-���-uo�r�V=9(����Yת��\I�����7�Xw�iHç���B�%U�#�5`����h�Tg�nnCUI��}����!��k�D܋h�;f�ĩ���n�TE��S $��T�,�v��ZP� �ew�ՐTI@��q��c����}8� �Ԝ -q��>)�s���At�I���/���\V�cb>��twb�3ǀJ�×K�ވ�����~�=��z�ً@�6���R�M�3,�{�ך.9�LL�:���)(8-�lҏ.E�� &x]!�%�o�	%�B�Ta[Y�UQ�k���ݿK��Ikq҄��i��5�7�S��-��s0$Vrx}��l]M��M��?���R�yL#ɐ���'5�!����ˀ)�m]֒��k�H����!PΥ��f�������t��G�u#��f����AW*lHSa�l�|&F�*;{ٌ�Z��Q=��g2	6�����f\0�I<[�8�FKd�w�-/Y�f�o�5꘏��US
E�؋�6��⢕K�t@U����
�i���`���F���4vc��ӟ�&�42)o�~����M�M�y�
�����	�ݸ�Iw�����@V�q�ū�؜�ʽ#�m�L�Q\L�J	3��gX�� ����_SV`����k�Z��G�4ǌe�-�Nf�Yԏ ��m���A���$2 (�Av*U:�����5�[�����b�i.���OٿN�b�nc�����,ɤ̰�h������QaӍ^�׵�&i$;N06�$+��S���N@��~��7�'��H��zʒ��H.kJ8}��cb�y�Bn�0��Lإ�]�}�B�g��9�5�>�d�c>��_�+��%���Upv�H�d

��g�]f���O��>����hTbMϘ>�wt���~�1��3����
O ]�c���.ӳ�Y�&"L�DD�:r҃��޳/nE��X��\��Η��׫-a���Pj_Cz]�����A`17��zy���V6�����˹��(P�e�Eg%����X� :c���R"ѫ�g�ˀY��ʇ�
�'֔��QxJI�X5�/�xT`9·�-���k��^���%X�2�0ȺV�ڞs�MM�>�N�8�S���m\����c0��j�^ZgH��S����� :�v��2V�*�Ct��R��Ȝ�>�������	������ͮ6��������#S�m�@�Q���͍}d�	ʀ[~^����[�y��KE$�/�`Q]=W�\ ^��$i��t)��(��W-}cL�z^��^��TӃ�ᵏW�~%��xO��9�d$�.�w\�95�ΕvD��vc��!pc����E��^У6X�T8���;�(p����v"���,����;����y=:K,��y��ao���u�[�F0DF�Y��Ib�OYp�ә@��&��{Y��n{��@������r_(bK�a�#�K����3��k�sJ�'5yp�p�Z��K4~�A~�f�P�*�p���/p:^c���H��a�#����I��_&�q�����b&����pd1��h�6L�٨�h��R�D��C�Ι<�-C��>ġR7�	�k��D�ؑݍ�>��,�q��	�5%X������V��[�D���͏]�(�
��f|0۴��ʔ��G��]��~J ݕ}O�d{��DtZ��1g�oN|Gf`��n+�W�HI�@"踕���gRᣂԮڗ���J��H ���tOE<�;ڽ�x�n�xI�<����R�mg�;�݈&Eٯ����G��8�3x�ɪ��<���@"���{UVf�%{�d:K���r�2���& W������t}�iAS���^P��3&�a��i��@MbHS���b��o�k`�kT����aD��2t����c�5�6��*�Ԍ^^M]pÐ����L�!�V�i�C�CB��q�+ڵ5�'�z3��7̥��}ul6�$wKd�i��J����>��V�W�����ed��3:�E���
" �F��)N�9�Ȁ��2d�zΤ�qIN�kd�P[�7ѡ���M��`B.D� �Y�%i�GU���<`N�V	i��/>��~2�;h�r��u�R�C�f�;=ɹ��zP�e����b].6#�d�d⇝ �vy|2_�N�\�R�+������A^eyy�ہD�^k�&��X�nq�[Y_c�=�¯K�0��iϥf��Y"����W���G�ߥ��z��ۃ��h$!1A����Ó��j�+���ӷ�8��yp�v��bk5U�A�Ǫ���_ճǩ 3:�}~܌�Ȥ87}4�<��ǳ�-��ݤW�ӱ��X��$xi��p��C]fj�u��L�Iko(�Z��*o{hT�<����{T�0����]5F6��T732�9�|ܳg��&�~�!��Sګ�{>���ى�<{Xȵ$u���@���\@;)4����AyI�ȴ��P@|��>���
�ܘ��Z L���m��/���� ��O·�+�Gq̓,4qPs�(\��J��@�镂%���i*�E3�s�6�7"՞�M�sZ�-1c���
��=��\�}�� ǩ�y�ڒf�Nt��99���u���-@[�}�H�^�\���Hl�b�_Q���������`LZ�&lJ�j&�$F�e$��h�_m3�]��h��^4ulS]GDX�t�"����D�6���ܒ,�몇��B�W�Ws����8�37x6v���)w?��������Tt�>��P�.s0IW�6�ó
�ᳬ>	v� �1�TY�{��^�j#�V�f})�3����E�(�^jz4����<���bB]Ѭ����u3�c��^��[}�/�λ����s��
8E���7��$$l�]~�i�|�8�t:��Sb����B��}�5��ͅ����l[c}�3��I�}�{���G���0+��k���'|�F(�U${l�
�U����t셣��?���NUi�ݘ��ߋ)6�g����u-�:W�/�W7L�Z�9ԡϓJ�8�L_��:H��@Q|�Y=�<����K�����J��Z��;����?�L� 	��p� �XI�˕�b��"ؓ{Og*�}�RK=�|p�$�����4;�ݣ8�keT��]ƻK���#O�-8+kTcq��Pj�D�]�E�Q<@G��v�k�`+#��T�ZIPW�y\�jo�d�)��0�n��Q����)ڊ���j1e �l���B�4�2�0&�*������=�a��=��j-¶й�!^$�l���o���C�.�]$�-󻊞�Ⱥw���4�H��Q�G�ʦ�u����������x�(�����r5e!oԛ��Q�[@���̠d��M�/��:��b���N!^��zăB
���W�R����c��<�͸ג�7�;M���{�~�	?2�(�J�f9:�)r���1��2��x�g.�AtS�4b���A%����AJg'v��y�4Y�������5����ɦ�unb��8\Sp�3ۨ\0�m��<�F^Kԍ�a�*��2��A,�c�G��u��!���C�[md��U>�7�A���*ZT� Tj���侗��6ی<��F�^��+��_��)b$�7@O���z
��؂1����}��,�r�N��Ug�zA�g�Scּ}�V1R�ۭ���9c ��&��S��6kf�,X��SKm� �â"�jS�6�9jL��vIuv�,%zs6#��F�2N�|���ׄ�����)�@�*T�4[��}t^���TG�w>5X\�66�l ��ѻ�# ���^�oKh^��}�#��wK��咬n\�8�UH]�W=Z��[pՑB�ୗ��.�QD�چjJ�ڙ껛�j�<���/���������*�a����d�?�[s-8[�%�P�%F{E�5�W��
�7=#XIg�F�=	����;>l9�a`o��<��x2.T�if�t�N'�P���.>���,��;W���!~<g�䂌��E�aQN�*U<��x��	��;��13tn�Í�N�e��=�%��OiՒ�Ѻ@�����]���e9�C�r y�#S�,���o�@;��(	׹�ۇc�
���W���"U�[�^d$U1�CS�S���Ш�$��^�J�i>N�O�>�*��(�0����0��~І�@�x*��H�B��U��xA夳."p��8I
�y���sl�[���N�O=W����Î�c�'���
y=u�;�2�����w���8��U
�ؼN_�$�} 1�ë���X�K���K���vi�F�� U����ϵ298��pw>�aʕ��n�*��(���pvK|���Q�{��5��F֋����9���z��"��|Y��!�j��\*�m`y���@�_c^��zvM��uu(�����WԪ�6K� $��+��=pї�8��~g�b)טBR���䝍g���i]��"*�r Dihȳ��r	W1r]`�F��������2@�q���ΐ	[�a��qoY~��G�_�.T�UD��5�'ٺ�ӋuK�O��*TJŐ/�qFT� �F�c#'��D#���z � ��(�ab,7����-lȾhQ�"q�8UjÌi*�Lލ)Q{_U� ��ˢ���X�PK�i!���?�B�2A������]!*�����b�%�LXYG #L��^�#�����Oi��'^�y�Ҷ�1.�j࡟S���0��3%pלּC��3��X��$o.²��RO܃;@*���4d_ճ(�q��T��~Ǳ�v�'�Q\���@щ����$Ƣ4��'���K�0K�,w>��&w��O��c`o�U
�h���2�n�3���^�GU΀��?��R�{���([��@7^1�1�8����%��#�k�y�zM���#?
ً�B�@��OW=����[B���g��� *�MY;�����f�D���#p� &d�û�&V���ĭ��y��'|S�س��dڃ��E�l�4��!K�	,D�&�_�w��_���"3�3J��|F)�6ԡ�t�!^���<�B�p��P���F�8W��:/�-^���L,�e�~V���/	��/�A�Qo��$�
7�/�-aW���\�
A�j���3"�!`O��<�pzвo�R�����
B�F�6K1����"6y93��ݶ������/q����p�s�\��'���s�o�4���P�L>�_KNu1�6pƌ����ϫ����%Dr�i��l���a�,'?��> ��#'�=��=�j�$9��AzgS�f:��L-�+��*e0{���mN�a�,E������T�R.A����a)=�qE���,�w�A��~��İ�������X��aX����T��d��2������}%�&��'b�6Kc��k}�U��m�ؤ��72r�G4�<P��ې��;�d����'�"�W-*�^��4�e��9XD�>�x׵�h�6#^��Z��9v����I�C��Zt(i���)t���^���M�<,�RPѩ�,��O.��tܚV{��X�vm��VW[U���,�ZB��=?�X�Q��e��޳��)`��Vt���Bs�zc)�f��Vҭ(��/���������Y�*-y(�K��Ҭr�=(qέ�Q�`��c�n�)��<�o����fr(�Ϯ��B�[-1������X�H-���\}o�m����k|���50ю2#"7?��/l��Dr#�v����m幃ɇb��M����t�2�r����:�֫�(��'�
|��5Y�*��zg�D�Е��H��g��^����`�u�&�ݙvD�}���,o%ѥ>�ޞ�24�	ʥ�b̏�u� 
��d����ŭ��s=�s�MA��~ޜ)ur�7B��x��g%a�G]�(���%�=<��3kE��\#|Pk���pf`�h��)�}]����L��5.v*ZBqr�k��UV���W �(yy�2j��;�h�_أV��}� �*�#+#�����a�6���ͦ/R�K?����pF�ҥ�g6�v���2��D��nL��ㆴ�ۃ �&<"π&;.��i�=5C�5����������>5�L� (���o��m��%�4ԛ��L��5"\͠���8j�O�ܷ��j��2�2!"���Կ��|J7A����^Y�b �O���q��U֙*&Z�r���~jZܐi"Â��ς��y��5f�CW�ῲr~O�aX�o��Eo�i���d�@0;���5��)���r�A"Zb�|j��s����Z$o<�������g��2�&x���C7�cb/؆�NeQ�r�Pu�ë���q2}��yF�@�@b�b�������K�>���Q�c~����%M\�O��c�\&�<Cn�0��̚���^j�Y�ׂY�8�q�1 �ٛ7E��;��$0��T^c��/m	�h@,����9�#66Ht��h+�qM$5�	�5d��L��M���Ǣ�6�tg+�
��%*qgBi�D�%���i��[}�/a�V2A���;4<�Ⴌ�D<�]k�� 	=�,���O!��»���M�Rh�{0�!��J�R���
�C���Vi�2���;sr�UidÙͦKe�=��
���\�0�{��y���3�1�em�<����_?{�A�MZ*y�7���V	V�	����Ċ	dOT���YLr�@�@'𲑣]���t!�O��b�b����4Iߢc�X��l���>R9뽩l�$�MTN".���*�H����*��ĵ$f	�=\�� ��{���t���a�c��� !Sm�TbuӲ)��v�I��w H�L��vɷ�������L�ԩ؅{>L1��0�n&*LFH���7�-f���,��{�U�d;n������N���u\�a6��D}�Mj3�����:y^t��Z�j�>K��ݐ��[���S�ɡ�:�V�3HdH��1�cY��C�� ���9�h��㕿b�]���<��P�:��jLϬ�;%�j����a���\S��˷���nί�T���o%Ӕ��'�%�i��DL�N�A��V��
�}��zmW� ��~���-fi�C>H���)���	��$ȷ��[9��`�� EU�'�H(�l�7�|��B�mHa��#��ƪ�q/濪6|_<4A��vl^�l RR8��n��߾fS����ES#9��ɷcCd�Z�Ue��g� _��w?׷
u$o30pЛ����>I�׵+��:�׹�P|��8~O�&��7߿��z�4��ƚ�u����;(�r&b�P@�D�Ih*���|m9��
��n��s#DU4���ec[�P���g��~�Sa���Z'x�0'�I�XN��+��Wٲ0���w�#�R�����'8�>n���©d�0�\
FM0N�
�i�*w0#��͆s��B�3o_RB�1i��m�
OXQ�JE����Mm�;%^�2�$EކJ����{U\�Va�*���h��7��h;cA�:V:��X�k�Ƹ� �|Ʒ�F��K��;exa�ϨN��)o]!��{�,qA�݊iI �b���. �̃wA؉��&s���o�@�_�H��7 Qj��CSC<�1��RL��h��`j����9F���A�xL��:�p[��<��:�����{�V�v��� /C:u#�hm3�g�X�x�=ƺ��(�Ʊ�����PD^q�w��1�Yb!QPcbo��U~�	C�=�>LoW�0����o8/S�puc�WZ��X���AȌ$32_�>}HN����<�i@��� u#Y���A*@�Z�U�M>�'s9� �^���!��ܰ^�RA�>UbnaR�#����ׄ��n�/�uY_�B��)\S���0�*Q"�������$�Otq��wY�[�K��Q��V&��%Y�_����TLA���0��VgF���S�>��z+�Е��2���`{;n�]Y�E��9�!��;(GԸ�J:�Ұ�TS�c8}v/2C�d����?�7>d�,x��9������~ku�,0H�V3I��F�\���w����4�fSz�k�<)5r��۲|�]$�\��O�\7�Ԏ��E*C
I�7P�J���/	�g&��m�R4~�A'� �nn(�CLH	c2K�G@�eH�d���<�����w��DSH���4�.Ŝ����"j�1��ݫf�6@ �ڂ�	�k�(�Y�`	t�H��Ú)����M�g���^�1�[+�+��1;��;o:�2���Z�K�z��d��+��rE
���z����9?&��d]�=��mw�Z��xS����tr�"�;���:�|��P!�g.$�`f�֓п��#a�Q !IN�%�_�����H˂��ӆ�qV!�z^����������԰���k/D*�g�廍�@�W�彁rIa�hh7�9D)���,����id��#��1o_!;	��A���1�\�3f.;Do�Rna]���ʐY�K1��^�����t[u��{����ԕ��P3�>${|h�d��וR$"�aHT!�;��}��J��b��*w���|��JЙ��u�u?�G�i������n��mېT���AR%�;�n�*��1���E]���BB@��%�x�ƭ+a���=;����#�z��k{>#�8`nB(�K0�C���b��0%_��l�RS�ū_Ȍl�ezRF�'�i�ٽV��S�L���֞��U��*�Ս��rz)�91�����`�_�u_XU�{�M7� pu������32oG`�/*|�{#-='�'Gu�1�ۊy�O���1�a����qWGz��M�?�7[���%�F��3\����3�{un�g�^x$X��c����;<髲ʷo�Тg-T4ѻ��lگA�7'��T�1�5}���V�*�����VPs�[�����6%��7�a�����B�.茛HH6g�a4�b� ��УSv{�����r�4�{ ������iR�뀠�����d�M�H��r	f}9A���rZ���{Q	�\7��6�.K�"���<*Nر�5��#�������qi��'&Ⱥ)�ϒ
o�?���2GS���3?�%�s_�B'Kf��
�9��7�򿔐!XҔ�;�:cZdU�Ic������,;�ƹT�>R��%�#���׾�.��~���&�ϖ��zOX��l����3�K� FY��V�뱦��)~9�m��e:��A��G���� ���]�+n����c���?����/�r�T-C�T�����ሯ�@��^fDyjn�ǝ}C��B�.*�>
��������4`��.@=`�p{�PL8�`Y��0s�.V8Pv�߻���֝�P��vn[�8���h�֚ŏhOD��Mw7���|�=C�ՙA�´�+�E|	��٭����4�I$�����iGp��<�۬mg]�v�m����ؚgE�Qۧ��0XC�;�{eR� *@��%��ý�J�;��U���������GS�QÁD;r�)�͓5E���lUCB�ɢW��a�`%�@l��^��i[�{m�8���{��>k��$�h���A��xN]�#r�밫�N��njB^�0^�!d������>|8#"��\�Ow�����V
�m��d�A�4s�:)m9���MB���T����R��Dx<�ʆX�t��a*�%���H96��\�f:8 <���0�ME�CAt\�{>O0�"�����O!*��e�.�k`�)��!��>���<���2'�<HDDVG^��×������q��Q�4���R[�-�o�3�ź�=ή�(�N$H|*����ߓ(�R�E4���z�1���e':8q��iWs�Uգ!,h_�#���@c�4�j3��0}�xR�y� �;!�3�?�Kyɔ�ӄ�l�.ک@�.l�*�S����>VLQ�hj�R�!Y���Y��c�򫵲���aI^z����|w�u���s �]>�-\���@ձŝ���Pƻ����^m�aF��x��U+��xe��Y���7j3�\4�mM�:< �}pg�3�(o�sJ(}o����%�j�njXK��d��������W	��
K̹���)�q�.^���]\�w;�=�C�������0c.䩧���)}��m���Ic�@^y=�ĩ]`�:���� W:ϋ˨$7�KrSE���I�]�}�Y~D�����7�&��.�,|��놲����g�%a���t������"^��"����T���n�T�����+�N	��4}�$�Y�_�,����Pz:s�s$7��Aj����ъ�����2�O`*������k��wþ�;��U(���W�)�� �B�*q����(��c�*���(%�N�Ih�ƥo���yTw't*���粒�nʡݤ�U�Wm�����+n����!�0�n��Y�|Ѽ���|�]�T�P�A�L�9�0�
p�FX���6���TQ�X�aj��c�C��x����T�Q�a�S���l� V��@T���i(�O�"���i���4S
���KT��=${�]�5���0����}2S$�i��!��Yg�����'bm�� ��V}�����&#���6��-<qrK
�M@�)ͼ�-�6�m�s�X����->Y/�<�IfU����d�чҪ}� A�cm[���\��`���G�P������$0Y� "l���@��Sю���wH�aT�\!.6���yr�����P�ي��������)(�'U��8�k5��.��&��-�^X�ҭ����m ���ӝ'R�e�%~����#���q��S2�q�R��Q]bDԞRm��������*�A��q�Ҍ���EZ&�!��%t�а���眿���,á~�����N�C;�GLq�,b�FAJ�o���f`F��U��(m9΍����,o̱���xj���A�~�!��ml���0� ʧw��Z�
,�Y�a����:m^�����Ǡ��ʅ���V�F���y
��l�|�!�8v�V,�e=%G$�)�[Sm�ů�icM
|5l�w1��29 f(�<!X�	RЇ"��&�����������5��>
�"kj|�k���~��l8s�YF��]pLp(����w�����z�~p���%
X���<�sx�x��ͦ��>mE��3���+��/f���5�Y�pnS4:={PηN�EK[V;�[ԓ�pU�Γ+�ݰU9U��&B*���չ�Z)q���T�/u4�x��r�l)�!3Bv�Ǭn��|��F����?i�L\g9��Ӥ:���,��N��:v�u3*���t�i�1�EqO��!��
�i�c���x�DYۨ�F|�8$x��V��g���ʇF�Л�r�Ss���ƅ�o�[M�V�b��b�2��Eq$s�+Z}j��G�*���6��0��C���i�i���Ove�I�;��0Z��A`lZ�1uTj�Cf������9E|H�>��q���7�G�ny�6�]��q�dm߾~�8�U�����蟏���VL��fԘ�ٟfL�&s:/�Z��(�e	T$v��t*A�Y��s�D5A=S�"+SV��ܞ���X.}db�׎A6�Z�9`���d���|�������#%o{sd*�%�?�rZ&f.�u�|8#l��C@�(��}р��_q7ZP�la�!D��1|���kENO'�([�O��er�&�WY(��#���Y�?���\G�W C�P�N��Q"��*�R}c3���TW�\-�?ge����s��0Я"HX�!}���C���3������ԟ7͞炥=�ި��J
O����I��35	P�Z���Yfr��\׾�M-��8qa��~��"�����~6>�4����ݾ�u}�c��FY��s8�F	C�%�:�\��w,�?X ���Yl%�Z)�J�"d�J�(u$���>$o��1��O�RG�m�jcϽ)��o@���/ȑ̤t&Nf,y��E%s�M�����>��\�?L����	��B�Z��i�XN��+m�᢯�o�N*�0Md�q_�6#��*Swe3���I���t���18#�lbc+W��iT��'a�˽[X���3H�}V���&9k}&�-��W۞�_��\�7�/�y�םl��u�4�H����@H]�[}eDݭ���'������@q�jj���M��po@�&�YT��w���cc�H���ܗ '�T�(%���5$Uc49ªs��ki�)��&?�m�U�1��)g--@�T�O�P�����$��y�	�~�%8�O����	�X3���o���Q�}����RB$1,)	����<�}� �n��E�?e�>7Xo�R�b������W��/n�<3N����O�R����v!.�b��?N흡v}��$��w���`�i��髥�� `
:�7]��S�fxnb��/v�}@��ֲ���"�m�(��\\?BN��裆-t���a����jOJ.�'�ag�]�P��)�e�T�J�_îl2��������v^T/p4Y�iDc ��*Vd'� ��W����;�4���╟�S�,3��W�6��y��R� �����7#�Pe�;6��E(����:K�buo�1@j�$S�A {�<XW�����z�v-��{�߃�#74��=$�� �p}j=nx��6��@~��MA��	��Y����8���,�#6A�k�OE�+B�4�=?k{�@�)6�-�BУ��ui���ަ��C����eV�	���p��y�ʹ���j�@��I� a�a���fD��Nt��
K�p�.�Vu��+�.���o�@]ҵ}Bw���Û��Ճ&i�nd����G���x*�l|V�,����A_�+<�M�{�"�_[���Xz�	�ڋ=7d��2��?BO�Fun 9���:�m��CO�n�.p�
'
Fk���"���+�i���Ӧur<u�zkY|"H��]*�j7�c��"���di١1GqUT�tsȵ+��Ϯm�L�\�3��׀��sO�@p'�ۍ�(B�"�A!Ȩݗ^,Ȇ�dÛF�Yf[ )P`B��}z���d�;�trF܌�c\X��ՙ�me�Y(�d��O;� 1�_S�[J_�>����si����ta�>��P�r�^W�&�;X%�Ŋ8oi�����V���R���b&�O^o��>�({�u�i�m*K5b塭���?G�������;���;��hz��D[�X9W�')�^��+�,ů���7axi9ROPMĦ����1�߮h_^��(F�ޒv�q:�6�]j˃�s�����@��$-,L�e@��~X݂2�g`����&;\f�ܐ����Ȓ�����G��ꋦ����7��$PA���2~����:�F�m0Ã�g�<`<=��c ��}-$.�P����ne��,�p��FC�>E�")�˴fiR�'A���L���ɳh93��%�~�y�[��wۭ�ާ9UC~�27G�3��+l��*��c1� X�&�?�d��q4!�q:s9*K�{�E!)����5�\5�s�g�t�	�t@S|���=D/~8�	�дҸ	��/Y\�	0�Q��2�AP]�A�Ȝ_w�I��ְp�������p\�zNי��!��zo�`# �����Ƕ������.˗�b���6c�2�;,�ay>E9���	�?M���Pڀ�B�f����K/9�%�[߬Q�&�7Y� ��0���#l�&L�����ƻ��)m{X�˳���]M�0�����Y!��>�ﲧp�q��eS&J}�N(� @�[be�ߧC�p��|��tL�Ԇts��[�c��!�S����,��~����Vڍzk;������  �@T�pW�.ۥ���4��S.��!%�S��z��a�!3��|��O|�pd�7����5i.Y�~oԏ�In�	{���
'N�!9E0n61�/��E�?�t�#1?dp�@��[�@� @�Y��K����sYB8�&?�xԱ��
(R���2Ȣ��8=�G�$.�vo"�[�&5��s��DU*�9���#r��[R�`T��`�xHB����{���LbE��P0�}o�m������Q����2�����0�axy�
���W�?�E
O���4�e Fv1o�7�An�.F{2��'���VP�_(�<�w��c���D
�T��5%[���
l�#S��"m�'�h�R������è��w�V��V����у�Ԙ�oW���I���뿤���A{U�괥,��k�Bf|C͋c,��,���啫+���Ku�%L�"9X��l������$ec�U��Њ� O���r��@���uu���܎3~���U5ϑ�.��:0��!��ִ��	W�=�^)P\���N8b�z��G������E���O��Y��	698%����#$TiD��Q9�S�4��T�Z/�9�Dkl����X�k�6�(uZJϒ�]K�d\�oVSx�t ZT^` �P2�'��#��1�����_���}��Kz-�$� �C<����}�2܄�#"�v������x�h¼nRÁ�S�e�� J��������P����cBU��]���J���LD+;(Mm`S+�ԐT��ll�<}���돈3��FMy~�Ɗ�4�w�j�
&4��ZًT�<�d��Q:<-��L�����]X��ღ2`>L�J*ǥ� qHN�ײy�H�J��^%���c�$�u��˖���I��H5������ AR��i�*���q�Y+0(�򔌻s�#S��s���[o��<��wx�9�4�;���t��H\�YL��Id߰��^��U���C����)��v����� ~�e���,��LaL%���𤽋��w������'���'c�O�'?<:CJ�ʛ�7��H�ǻ�6�B�Q���������m`kO�ܨ-�}��!3j���D�ʺ'���	?Y��nWSR�'�ݣ`\"�ƻ���D˹�,�zͱQ��w4ˋ�?{0�]��!_Z'ί*����)I���c�v ب1��}&Ls�IC��$/�:��2��|C?��4�^�^�s��{gg��{���~0�V�%�"o�0��؆F"1�J��ѱ�$�4�zKV�
���O)�#vB��V�2cd�<��F��ǹWX�k��B.��^^M�=,F�]k�t"��}�*�C�aﵥ":P��{�S-��t��XN=']�9���/�j��͠N�+h5��9�㚟^ڥԨ����>������=ؽ\T�縆qd[	N5|���,��dz�N�k��0��J8"�.VK��:Ω�tެ�"ל�<�ߦ�e�ɭ���<�ʇ���F�dH�+BLU��ҧ?��nM:��}fH��?b��DsY�ӼW��0�@S߅n��ͦv�j����+����%YȂ�9�k��+�)N���S��ɲ�N�5o�E�	8Eނ v'��^��7��_��#�nwVF*=^2o�]H���3�j Fdan@�%��	�>)��?�r㿔-�q#�Kw5�s�lq�6>��̉�|'�iz�@��&�5e���y~����^ a행�hۼ�����AmH��Gi��q1ֹ��#�asg��M�nף`@7�q��7�oL��`}�ȃ���g��)g#!}d�*,��B� 	8���%+�3�rp�+(�"���|���׊k��:�E2���e�i����h޹�jj���b�w�"�j�P6����;��i���cf����1�gNH��e!MH�6�_��!���?��T�Z45�ɨ0�&i6����@C�M��Q���A9N��e����:��AZG&p��sy;3��x�k�H*<�{LSr~��mm��z�����Qzd�x7��������|��'T���څ;E��K�:�I� �� <B�1��X@�I����v�������g���$�d���O��Y���S���c�����*�^F�%H0 y�XE����!|�gn.	~0r�m4����>gǪ힍yw+�l��y����]�d!\�G��-Ѳ�}�r6�sl�}���IXc�y:�`N ���!Fb=��=�Y�޻�x�x�΅Z`h��W����T�4=J/���Ogf�ʹ^��:�1���i<��է���ƭܗ��1d�&�7�o�ր<�^c-7���;���̈́�-�f�G,7�<߈K��J
1Ȥ%G�{Yhh64.���yR�u�a�0a��
S�;:��r�I�P`���7V�Æw�B�EԭnK�kx�tI
��#�;������uZ�9<�s�Y�U�u�B:�B<x����9� T/���~oX���h�>���=}�}�$=�0M�N�Z�g��}���)Sj=8K��M#�E�O��2�谆qp.d�-7�u|q��	k��Sy���#�g�(;D�ǗHLl�Y��"���ݷ���:i*�5wz�N1V��
��#��LV������'s�D�G	��w������^��1b���W����M�M���'�EEų�sh�B��T�H#�4$ë �@������j�;��\2'¨��!��W��2}	)��5;`4�T���`�I�¶���Wk�?F�-D9H�je�?�Ƣ�BE����[���~�l�t8Q�kCώ��ʶ���1'������?��IeO��G1Z�_nb�h�lx|�H��=�5��h��QX�բ��~3uI}꓇��
l���
�Po�%�� :SbΒ��o�6�P�s�gf�	{�׋m I����Q^�Tr]��9�ݜf��Q	��~"�.�{/C޸s�89��D(5f�|e�B��XIn�������Әp�����r~�mQOdX ��<lD�n}�O�0�V��EK�^��"�U&��������ۥ�.l�t��؉�A�)Ex��̠Ky���6L���'�~�%bԊ����ذ?�"޵�Z���xe|G*4dʋ`�����=���tc��G�W�_3��%�ڣU��Ŋ�^0\u��c�b���է-�c��z�i=ٜ�>J��:���)<;�@{������=�O�A��%ᔽ`���}��$��)�*�Z��k��:TP�ɖ�LPs�(����`�T�T�sz��M��r��7�!�]�3�1��%'�U�A�Rj:n�>u.Z�kx���zR�j�V�E�443�vA!MƄ�ݗ�s�Ve�ˬ�>�=�^h �_�����0mm�:#�B��7.>���x3a� ��^��vn��H��T�6�mD$=�7p�����
��6D���f��\�n~Ж���o�;K� ��ь�Ȑ:�_�aYY�>��B�3t�UX���#�O� �5����oz
3�F> �Ʀ�r��u��-tw庣gnc��$�1����	�$-I0\�U��$�n�>.p¸-��b��75�K�m����I+#KW�/�TҼV�x�r%�|��#+YA�rV�ܗܴ3,U_ �����*��K^�����()T3�x�YY�2QM�f@���Qn��&��� �� �opS��a�ڀ��)�T������� )�3�~����Q.u�~Ca���Qd��=#X��A�In] ���7�L	q��ߦ���<��ko"P�g�ݘ��~?c����m�3}�v�(��|]��=A�X�l��s�+$�l@.��|s� ��_��E��kڳs�7W�k�x`y�S-W�N0�=J�o�f$���\�k0�·�����������s�7Ҷ�Jnj�G���f�{he����L�@�i`���U[�іC����:�EA;;��C[�W��� ��z�)@�-tB�`V���OM3L��>T �z��=�GRmP��v�h�G<�ծ��3l/Khܢ`#�P%	�"��9[��d�5J�j�
�����������b�ˏX}�e/�C�QM�@�G݁���T��f1�EK���I�)����:����.��+:������G���O���K��R��9��ظ�w���!jn"�����qB�,ŋF+Tyo��f�v���	��=&����Y$&al���2�^�;ҙ>ڱ"�K�t6[���bo<>�?ȓZ����cA2wa�F�A���h���&�iJ�5��g��Q/����P(7���
�h
V혥W�p,M�#�/��t��/�j	3"A�W��� ��r P �^��;=���TN�*4k�=�"��F���vw�
e>n�\�m�"��'"?�Nk�AښO�g0�9��b��o�в��8�q��qW�IMj�j&�<F���"�j�#w��}��Ðew�{*���0*f�/�A���p�~�H����������6�Н�.�X~Aܵ���I`_6�'�󍛂�8e�b�P�.-J���!DJ��j="�O2V|;��U�X������$��	,����1|/�m0ԙ |Ch���[�MO��(H]�<�o�|�J�%�G��pk�`������{�zT��4M��(\��jv�y���ڦɺ{��|�rl�5C�(���Y��J��xٴ���x�������Tl��80 �$v�@x06hZ,%�{�	Crb�K���_�K���p�I��o*�K"�V�����:�p{զMN���C�S�$�o4���uZq�t�c�&ԁ9���(�[B<ʞA+��[=�Lv<<�[䥘q]`B�Z�޼'i)^أZB����;���l�vpA�%CH�{i-.�][�>!I��c�����[����5>�?9�6甸q�^%�2匷7�X�F(+ ��)��Ѝ����E�5�Od��i[%e�3�k���7ܞT���W�L�Ry�J �:�k�~s;��ai���#�r�4l������#�}�m3����d.V|̢3��9ڴ�;�:UL�o�%PW�ɸ2G�B�.3�7���8��;_�̀�6V:�����ɂ�?Yٵ;�v`���~ِ��M�bi���O�h1_M�j)�"w/����v1;��q\�lϋ�KM�`��f����s�u^ST�"��ds���ˉ��՝0�jL��nIv�2./����Eȴd�v��i١@ ��g����|ݙ�@.��)�(IE��}�w��s������{Og�eɧ�S�u�HS�T#��r�Ŀ��$ќ�ѡ����x��*��8hTjk�<���:yƧ;�u��a%73��"l5z�@�5��x�A�ٓB�"-�Zw���&X���	�L�Z��0�M�f�/�Sŷk�E��	+3��)xߓh��]�~)Iz�Dռ��7�<��.����� G�>�:^��t@���u����,_{�w,��j�M�r� ̟���ApĨK��K\�D�UxUq��=8�w ��ڢ�݇�-K��,G`i9�*�n�?�������V�n�&l{O���~��;�U��-���:>�U0:@���<��ܿW�/���o����N)6߿��5W���.�o�?�)T2����]��y�F�x���C!MlK���ls[C
�?U0�`�t��ŦǗ�Vÿ�vA{-��3��i�ŚSp�k��D1D����u��`��8>K*h�ޱ��r�xl钚�eDB�R�
!f̿�R,�0<$�wdh�����J@~��m�?G��z`����vkz��F��*��e�M��F�{�^ʔ�C�@�t/�qCeax;"�5����`��:�w�j;��	e*�0ɴ݄�9H7�$|~x��k_�ᬦ����˴!7�rna����X G&�R��͑�����ӳ/�f��)J"k��SO�����L���h;W��$�ď >Li�"�61bo�h5�[����KA��uz�h�ֈQ؂�fL��Ψ���������B�ث�}v2+��Y�p������[*�%����{��������6;�c�

JI��`�YG-�#X�>��v���[�H$���u� �+`U1����K��~������F9������K$I�$uQa݊�>W�z�"m�a��#?J[��v�[Oo��ٜYE����A����U��j�޶�@ŵ�{*�^�ds��9���f@e�&T.X;\�H�*m��hҵ3��|�2����>@pz'����Z�0R�E�	%`�e���՜�
0x��V$��|�O�[D<߻�0�jE�7a�'�D�-�������О�5jrD���V�a�H?V��e��J�Nu>�U�#s{���1��T����m{4�J�����7������gRk� ����F��9�*g*P�v����t�-�mY�@d�u[�Fh�����TƟ���
�9���2�Y�AY��|�\�-�ȀCU�I{��h��m�������yjhoX*�r4e�#(��@a%3�����+怼�¦8���FOh�<ykѢ���&TϹ؛�x~����T�������+��v�#`�Ѣ�n*�ֹ�Ї�����E?b��q��V����T{-A�O���Zd<������Z�Z�^����[�^7�+�����K��{��i
g����ynj�P0� �c�ZX�s�Yjh�PA��[�Ϯ�9�8?�$t���\J�.}f���}��j��h>����3�X�"�jhm����5�(�މ�gw�\�В����kr��[�B#v�BbD�Dr�E������Gn%�臌�k�@��x��Y&��?
 94~3�AYS�%4�U(�S�ӥ]P�� 5��!���M��%Kk<� 
C��>�Uˌ""�,>o�c������K�9���\�Jys\�`+����TǇ[V�'4�
kT�e���B�=��G�d�IN��F�FJ��4�ul$��G��g��m�.��.<�f�����<�/cg�:����-?t���{�b�<�u�Η�6��[]p!�Ūz�AY�InkF��m�4q���im��V�V�"�f���f��:)�@�wm��� ��.��+�;W8�K��H}��0����XvRS��{$�����/e�9��s�Ul��s��q�����"����v(ô���N��f�l��:��b|������=b�J�;��j�/��N�%Z�h1�։��!�i�cW�8*=Z�)��a�%u;5A����-��ۻ�b����B{zF"���X�]����ʭi8�KHY{l�)i�d�\�y}���BT7%Z\/�R�CE�g'�*c�Tv�¥5�=�n������T{l�����
��{�;)�0�&�Dr������P,@�g|�9��r�j��dGѰ ��3�ki����Ս���
6���2���`��K�h���kxxF�/�.��d�J�A��T�ǳ�?hZϩ
2(��/Cq̷X�D9�\2F�8��2�;��3��ٓ8S��㬵-�Fc�:���N�HeP��]۳�<�I1��e�a�P�xk�Q�K����8�Ej�����5�
~�J�|4{� cHҗ��7^ss�`�����k�����x<P�����t�(�e{T�K�n�&����W�=���Fe���>�B=���^�Aek/H-j)4A\�=�Ǖ�q�9��z��(����\��q��N�hX/ḕ2��H&��Bal%hU�����\+	�Ԑ?�>%\E+̰)rM�����J�F%Ш�8^�S�����X��	�H]��0?���|l�I��E��O,P��C���u�5���]��3vR���O�h�nC)G1`\-XNe}�7EBoJ}��0���#��h&���A���VVs^�{�$�B�j���	��[�0���d����4t1e�c�SꕅJ���+7g��h�<�� јJ���}{�۹�1:M�%k3�ݪ���i�̮?N��P������Yjx9#z��i���3������;�S�l�i@(���� oM�+�������p�P^ӵ�_��Uba�q��''�m�=��--� :�����{�Ԏ���1�5�r�)�q�	���|�N�z[b��p$��B�����kAk�nl�H�e!l.�A�I�4�{�CR[�蟈���L��zV�=l'9�<�ǡh�͖���{�\��iЈ��	˽�S�/Ώ������fS�0 ��B�ږ��6�D ����pO��w�I@fB��^��v�8�{�?!e ���Ā�)+	� [Q�#+�kM|�$�8�e�]3O��d,�}�?z�w�_&��5�(�����A[f!P���	n���o������!�#ru)�(�c<V4���e�����3n�;�KH��p�훗h$h	�A�r��%���C�h˔�{Z�8o��[��%�D%ށ�7M}ۼz��]4m�cL�7v�->c�H���7SNKO��q�;�N���}>Ȏo�D��+D��A4�!�%q�J8-��e��0!}��~�)�:�ۍ:���?%�w�$6��W��˞��
���>x���C����Grla��݃�4�b���1r�0�N��+V�u$f�qs���n\'/�m��Zs@\�q�<�^#��"�u�;�){y����(oLDR������0"G��>��V��ܻJR��c��|��M��'DA�)�Nt�$���Ze���;$l�'G��i�,��3g4Z�^�l]Zv[21<���?�z�{��f쌆��a3�J,�!q�눍�b�y~��R웹(���L�*�{n ��"�r��8��R!b$q��2���ŷ��c�}6 	زpA��|<Z�Z��3�w0�����L Nv?��5��"���G���k��Y����|jW�¹	+Y t(z�(�RKC��B N�xέ#��AFH@��;&���a�B��� �9x�uǡ�ֻ�$�iR'����7G��6����?<qu�l�["9���Qߩ�c��6os��xP�*�%}�Wȉ�x?2�@z�,�Ǌ�lKSYL���[c �����;�.L�[�ok�&*�E^�e��� ���pR�on�J�6.Y�t�D���Ѝ�$���\����ʦ����H�ZF�4bIB�rN�5��-3�P�I��EX~�^r��B�1]!�b��@F��J~�_���UX=;PCqX�jL��f�dE����HM��#�0B���p^���C
�6f�`�Q�&c�n,�C&�!�4&$5��R�)����<�'�G��
�M�hߐ6i�ٯ!on�N��܇l؝+�-Y3jC����x\�Rw<yʛ~_2�1V���~�\��b�F��@�?x�k|"�V�Jo��0Rȟ�������#DD���HE�P׹}��r��-�	ь R����;�/f�wD�㔺� LP��SƩ�W��M3Mo���
ۛL�'|9VV��m�[�&�@$�һ�:Q�h^�]���I�����D�v���Ӯj�Q�j���1)���.n�Zdl'���B��j�UǸ�%�w�/���t�gH�<?�K}�\wl+�M���h�Ւ�e���3���A�G�DE�b:/0?�
�FF�u�>Ѫ_�
��_�k�M4�!u�)��<�/��/w���%-�{��ɪ��ͣ���sQ��	4���"!��Q2�����ngdЮ��{D�0�%9l2ޥU�' ��JO��/FH��Yl��B�$ΏܻzE*����oĉ�E�*q���:6��g �k}� c(#����� �P�f��d��k�Gw��-G/-�9��QUVt?|��޾��x�B�kש��� ��f��
�]�"��u�� s�a���iũ�˽i�Z�q��0!�ǒ�}j���NXD��gb���®F�
ׁ	����\����9�A�����B:�}7����Ǫz�� ��lR:W�NP�������ko�YO��ZT�#hz\����N^�L�.c0|Ja�P�)v�xQ�u����E��Wq*�F(�1�]tV�o��(�6:��|�ܬR��M!��DO`k�kqu�@�_�R?��B�c��I9]G3���>�ԛ�p���s=�ș�������o;\��W�k�8�8����%���v{�DF��?u����C��|uS�JڙH�i�� ��@���{z������+��Wϡ:�
'��� �FG���N0��VYb��_"�������y5�w$���UQ=�A���HZx��߭U�S��Y��N�
OmT��V�B'�2 F�t+)]]W�Iw��>:��ANy �܉��C=cWJ-޷�����ji��������l�Ii����jK�a�$��߱�0f͋wZ͹�^l��������.�� N�nB��Z�=8c̋�A�/+`f�ON7��$7*3*���O锺�G:T_B'ji���v
�y��� ��/�6T3�h��x�vC+4"��F��_��Fș9��E�_2m��*�D@����BQ(̤��z��]r=��W@X� F��N��[˥��N
�p^���̵"�����P��h��o~��T�̹�*`7��6�J�(�B�v�`_������!,*iڼ�_M&IB���������4g�~A"�W��@]Q�5[�����<0����ŵX6!`Y��p 7Rkn���	Ű�����ݓ�W��ˋ.߆'��f3� �'�B{�Bl��(�*F�c�7k�{F����������_���{N�Mt
�'���>2�b��V�ڔ�| �6�	,'�W����xr^�q�Y ����(-��#�� /�������N�+�7R�ku�Ld�Y����������F��M�l�6ZT���?M<���ײ8--�f0!3��_�N-��0�0�9�ů'_��w���A
�/R:2���/����
5�5Y�x���E/���:y,�Y�2r�y|���
�u�Z��B�=b��Ǘŀ�z�_��X�ǝ$�����Ԑ<�/�J�o��ž���1lT��/��0c�k~&J���̙�yX�-Z�l�i���c����d�?�6����G[�b�Y�/���� QUt����)��@��ы�C�c��l� 扎�@w�f�'Y�TY���Qr�d�p�ӈP��=����<ꩋ~�DM���iR�ۧ�=������>Y�A��S��D������:W��/�.�����T���
8I�K0w�$J��g���wz@w��^���iѠ�d����YX��5*�#��u����5O�dU�iM�}mb��� ?�R�u
�q����A��#]�-"��jM�>~4;�9Q�����,_F�U��VU6acM���G�7IH�<@�G+:�2FK�E�'n���E�SY����Y�a���X%�:�ϖʼ�e?���s��K�)��G�n��N���917����z���6Ja[�ܦT7%7�����O��<�{�S��)�Ǔ'b���=�L�M�	8D��Կ��.R����#�e��`�K$�W��1%��~@NO��MQ���b�n<vo��َ�5 a/��W��¡��a�t�*�����ǯ���1���$Y��yc:b�>j�+���8��<�t#��#�'!x���! �*\.��O���u��(T�K�Ր�PQ�����5Z'�0p*Osq�s)�3�W��l˱�~;�%JRa��e[�[ʾy�
�@��������"g8��YK�2g�Y�tsN�C_1�ք�C�0�Z�/����D{I/|��D���q�"ɼ��j���ʺ~S��B��A�^����ȃ�a�hcU�tV��>f���M�7͡�T]��� ������>rh����{z��8�wȰ <���y��q��Ti�ƌ�7�uDWt2o�#8X�l!iQ��M������r���Á��*=��]�iׂ��⭋<�8����=� ���&���Z�B@�{���8f4��;l�kƩʡpo��#��Aj4zxO�ˏ�3k��UӀ�Y��WYm�.[��F�SK�V��{�ab��XD��Ȫ��>�8�Վ6�
*\ZѪ��L��҇<^k9'�Xt�����x� J��ΏRD�=foe*��7�6�A��Z5����|�[�����P�$���o�ښP��������l��{�c�(��)n�x�#|,��������>���� �=yĦJ�Fs+c1��mR�"��;�>-�䎗�0�����N�ĝ�o���*s�as��0����`�P�Dct/�����Ug�a�D3"�}��D�%��qF���ϡ�'Jz����묶l���:��(���'��y��%A�^�* �� L{�X6r�씃�d��D�N;�A
Yai.�'	���(ݷx�Z%2�O6�¥eRb���b�Is!��O�w�%[���tY(bW[� �$�g���ZZ[ad
��/��b7`��q��t��An���H�[U��8.*���c�޹E1��8�Ӊ̷��!~����m�v�QM=��-(��W�ǯm���Z���N\�I[t� ��R��E�2�;7���* cK�)��C	�V�A�ޗ��(:�W`V����!��4�̧z���O��
�G���I���LN^�&�K��2��V9N�Lj�~$�>��ѵ�0��<�O������v`C��=�9��Q�,r덓Uur�BȀܾ�.W1v� ��j�$���1�A��3���Q�H�=d�C3D*�۫,>���A���g���J��2�64�l��]ߦ�#\Ws�V�C��p��"L���A ����E�%*�8Z���oX^۱MRW����0�I!/�[sbhF�8�C��`"��&I3Ey�`�����׭�fo9�4�=b�c��"�E0��ب2 �h̯h�����:��&��z�� <KF���5�z�of����D~���l� �'sĐO��Y��#	�W��
�匭�A���ec m�E�r���d��׏�<���G�v�oR�5�2���[��*���W �BT��LF�?�0O�bP�T=���QR��6�ӒGӾ])�i������qxKؕ)�t�d�ZMޔP����EX����/F$���w�@E^ 7fle���@��'�M��3���ɶ���Pw1v���g}��,I�p2H�,y"%��G�i�22�"bK���Ngx�vq]����ӄzp��LZx�칠|q�I������5w9�̺flVgw$��2{K�Q�҈�v���}v������k�,��7cw1��j���!�1T�9�Q)��^o��P�Ȕh)�uZ�g)h�P�G�9vA���K�@�Aܹ~K]D�Zz�6U��M��Qves�a-ו�a�k�:U�ƭ�}�[�.7�|_kOK#�����=���-x�t�wZ'�4�)�d}k��+r�%��k��oܜ��!v��Ih��5�9�̒����.�Z�OSyS�Z��8��*����~��' ��h|�	�ڄ��a���e��	ԭ�U��3\�����
���d�>��*��DeNvԇ�����JÓE�����'`�c�dIȻ|�5\,�>aO0�27a�G.���m�q��uPH&|?
��l���J�r��v��c�%�{�l�����c��6w���7�r���Lla��jW�\-$�!af
|^��y�d���ܲ-g�d�/tm����N���۴&c�&NЩ�;�
�	�;-	p7�m���U��H�����'wu-Fx���\v��5���n�b�~F�J����,v����/[${C���`ne̥OiԊ��aj+۩}0�w��>9q,�JO�kν�6S�R2q�������:��g��s<J�g����5.p�H�Th���o� �oV�ʰ����M\C�L�����0��K|�
Fj�<\�q簸j� z٦~Mġ]�dI�S�Xְ"�8�r���EAɧL�_��9����Q��~�)���_�sId&$�D)]�=�E$:ېK��$>���]��xDxkf`0������c2~��Z E���3+����;���2~�m��O�����k�xiR?z�� ԁ�~���(H��n�M���+ny&Pc19���Mָ����_�`��<g�?�9cX@��}e���\4��fG���`�%ڂZ���N�B��
��ԭ�G��Y�_I�hw�ߢ��|��C����,�Ia{��ˍA��g�\�lfr��L����#㪞{ }��F�$�sővc�UL����6�~�����|3 �J�R%P l��� q���}ɕ�,lJ���1;��9t�D6�w�l%���툅#�@�\T�&!9�H�������J|�-�����$P���.Y|��%*�G�/����֖�d�s%����{�
�qXFd��@���
wI�f��-u��c��~q�L�g�j���~�;%����a�����Hrl�"�c���>�u:�)4 ��e���؊_�i�h�M1���H��/͛�g	�<��z	 �I��"9�	33_�	t���[��B��PxZ�:�/O	l�@�i_�u�;�:��Q�(,�;�� \��w{Oh���<-"���~���d�AZ��rM҆/���M�}kX�2'�>���Q�e@��iȀ�ƛ3Ni�hq|��N� *���4��iz%цI���1A�,��~��\Q"�� �$X���F�e��عz�z�^�҈�'�%	�����S�ņx~!&�A�"��
L�d�w�7�x��`�q�܇�,�+�l�~��Qbɤ�gri����Q����~(�өWnN�*M����Gt���ގ���$�Ƭ����7݀�/WL���>g�C��4���X33��!��rkM#U���9�����Х�|w3��o*�#��L��	�����!.&�""6��\�]��ܱl����!b��������������7m�q�������5O ��Pt*Y_��|�.GH���Z������"#�P!~���5!!P�p�Gm��K����,���\Ԉc*�WWG�J����K�Jw�V-�ay���>=R����]*�d�?�p3�X�#ߋVŢJ���D7��G��+�pU�r�����;��P�2R�5��7�NrI-��8��!Яb3�&��ǘo�t���:���&n�d�])���\nX=F�5cT�3� �Vv�hiM�ZNO����Q�A,϶�:����kR�� L!�E@�����$�\��Q�f*N��jF������-�/��/B�A+���s�rv���:����}V�ՂA히yL�/�U���Puh�~tA����epj��t�[�0Q�	�_�;��Ɔ�M൚
�k���cs�fM)��X�|�l�ì���s����H�8�ݍ��
{�M�Ns��_r�~�����t6�iծ��;p� ��H;0^�\���R~�[�l�?�i��;�2��,�8����`eQ�K�گ(�-7��uHWu㛭2�������/CU ��9<m=��`��5%��u��w$Y�@ܙV�u��������&��b$�ݹ���;%si�qy{��U��k��3��7���M�)[cuNz���y�G�EA��$M�(qı���:1TBI�V�I���`z� 	�~*N|]��n�D{f\���4hR�O�|�g0Z]���	ڪ��_�CM��8��5�d���D�`7n"Z�z3�C:L�<�ܱ�T>����F� �;������y����n����7���u��k0�����1��d�Y�!�*�E�)i�=�;o(��7�T�޽Q����|M�����V��a�.Z�vz�Ҽ��l��@2~@���Y[�a��M���d��#��@aL����R���iB�bL�+��A��VV��,ws��\v��&�~�:<�/#�&Oma��D�V/.��T�U=�>�c��0H�i.��o�&3��nߋ��J�#p&
˷��-�Ŵ+��ƞx3���Oԗ�;�����Yp�F�����0[2C���؃�{68�V�e�"����
&��P���?�i��n��
ҋ46�
X���u��~��v(1�5#��L�sQ����3`i���V���Ax}V��ݒ����'�RK�� �C������c�-<�xr������f��)z�DnЫ�J��U�Y���ݠ6�����Nv/E���;H�b��-�����XES��tԑ�� Mi������'@j6<�Ҳ�6�v��:�4��,=ƒ/2"&��_ G�(JK�Lvś� �W�@�3��~1�D�t[�h�m4P��d3�ě_Г��
�qOhW�£���P�mR���A�����p��	��LO?pKbl���Al���	�i�*�{�+ʄ�Θi�Œ]HU�����;�Χ��6v^���.\�gO@���o?������`Z�u�|\���Z�E�@2 �ժ�?��p�5N�M�]�r����i
�hV�$��H}(�7�]s��K�Ѓ�L*�:�r�g����mt�DO^2�����X��k�1�eo��󰁏����#��Μ�Mpڵ!Ρ���$��vd>u�ӿ���lN9їt��߰��|2�ڟ�25'f-w���[K�����.Y�ҡݝ��kK���K����NV�&]{���X�G}Kԝ������cƢ؍��v�8D0W}���I��hˬ����>�xM�l�9��59?��ɲ����U@l��J�r
��Mg�ׄ��@nV]�9��G��@XB�ea�����{�-@l�T�Y[!u�5��&��]2�n[jL%�Ocq��	R��2�`,��]��D����qi�B�ѽ2����y:U�+���u�i�l��a�m��l�j�=C��K��+h�n��ؒ��{=L��t���\�G�2<[�R\L��j![�N�U��	���멋�^Zr����V8n�S"����p�SI��7��S��в��)����q0�ߣ�^��.�n'��l��,�������)��C�5����+�"lN�i ���p�ĕ���I�!MYZo�Rg�a�ku���nPr;d#N���k&J�j�80�tt�D�Z���szb�7��m�%�{��IB�Λ�3��KMo~[Hë2��V�~oc^]|t&?8]�7��F��@s�k��9��k�}�Υ���|��"���{#*jW�&|�?��-��*��.c��B9�����~'�U������=@�ϋ}֌�Ce��ᬜޣ,��(,}��2�ѽ��#��YX���f����J�[ ��{����0��w�9���۫T��#��i��X�Y�JSW�v���h*����wo����hm���/��:�
���98I��kj��T��R�!-M�o��^s����p�|�T�Ѕt���Ǚ����m�|���(�ߝv�[�&i�5���@�ď�|�l�L�X�QUv{(G	�Z���݈�q>�r�u�D�&A��JSu쐕���1�A��.}"��,��RL Jmځ"����q}�.��������U�k*\?�_�`�n_�$N��{��D��ћ��+�D[��ls����v&:계�0K�Xc�����e3ʾ��꿾�$
딟�x�[�Ik"��6ߛm���H]�7~#�����I��O6N�!Q5���}'9����,����9�Y�ȍA�A���F�B܍@�DĦ3�1RX	��OST8�t��%�=!J�.���1��2�M�,�N�h&����u�ej3���DWV.0�ĒrI^��@X;V]�X���{%(YD��@V�@}�o��&����Z�^G�'e�ȩ��VY%�I0���W����{S)�W5.�r�ǅLE����A�ֲU����G֊yB�i���@����2")<n�86]F����@{;�3d�5X����_2�l���S!��]��*.�4�4|�M�4�ȴz5��dJ�����2���*���#v[�v�����%�e�� �K�rN���h{PS~��<9�;��o���O�1*������ܵ.}�D�iݺc07Ā�MK��ç�o,Zߺ*B���Q����g���5�a���~�R�馦;��F���$%���T�F;��P�uxڐ���ł�V���Zb�Rս�W���6#�o�U�yTnX��_g����]�a4�s�E�JF�Lb�4�<o�i˧#JP%xM�~�g6�F ����}>%��gLn#K��ˏ�g���r"ཨ���G����@�JY$�>��+��}[>Dc�HOG7Q�Ȍ%�T�:��Fi�ݮC21�tA�<Hj�0ʲ4��mY(�I��{��"����p��J�����Ǘí�X�vՏLm�kl^��b�����tŷ�߃�Q�?��0�Q����n�+b2=��|&���M7�P����G���icnsl��`j�s�=�e�x��5����M�%�1h/��݂�[Z��i�!0�	��i �W7��m��\ijD��|���S�MG�S�k�1�x*��%dm�#&n90��T����Ѻ�*�4����,�E�g��zC?Z5�'a�P!�JY��OFPZ���.{��1�k��:X<���������6C�(��_��� �$�N!Ys��o�+D@J6��8��U&�խ4���C|�5�C��fS�d���  	EiWx7���=8(�,5�'�&��
/��]�1���X��&>���m�`�Д~����]�E��QVp��V;����x�r�Z�8UC_�A�%��������K��I��&
û�r�[�x��J���B#L����Z���'�������c�g�z�CV~��,�)��:$$S��L5��
�xhv�/��̈���@�=$�F���{��g�Tl�m
�u@�W_�3-Pf�ROS������?����Ɋ;�<��x�S쬫g�~�:38R��czB�Z��,:������ѡD!����¯
'��q�@"9]u�ek8m��"���KA��QH\>Ī�m���>�n���3���&s�� ��z��&�T���L���Q��#���g;�c�	���3��8ݫ|V"+O����nd�۠58y�<Y�)]F9h��J�>1�ؒ��k�w���vm}.�W���-A�ZtPO��ܹ8Gv�� ��,wx�\�x^�W&�X ����g0~���gOW�s�*@�[���2%Mv�4|���`[Q���$�DH},	����Cv�j�k��
�.��r���Fm�z[BB
i�h��L(�A�L��NC���|�v^s&�!�G�&j�>�Ku*u�U�fj#�b�Z��Fm�3�`gނc�p̷��M&�����j��ĳ���u�8'��ͥ�W{IO��@�sK&֭�ܘ���dVq���<b��tO��v}�okB���Fm�5oe��^*?�p+�'@�%14��Y�w���Do��8Q��g�o�&+�l-n��9m���������:�\����iW���Z���ٜ8M��C	^uͦ&\�`� @�|�kd��5�K��k��r����AV{z�G"�4@Qn!Ӌ{?���_�_����!��jË�u;=}�
����W�Ǒ��NT!r~-L#������1�5���s����rH��M�=&6�Ήs&.�6E�]rA�E��;�ss����B�4�Թ���o�������uŇ�Һ1j/1@pU �Г � �,��9�_?@���3�#wnf`��Z
�$ �;�99�W2�ږ?���HI����*�%m�����W��D�M�9�8���7?�o�p㿍��*���V��pc/�,z��+o=kp5Iu���*�b��l��V��$[��	����i�3��	])r)�, g��`��y/'��ȷ�!n�O�N��I]ػ�ڭh5��!��{�򕙞�����$�8'�j�@���"	��7��&�̴���{Q���̓��p�p�7���
����N�	I��X�&�ّ�����US$o�0���p�$�LO&Ap2��Q���������D�j��k6'~�=�^�r�3�i՟�3*��e��b?[!�@��;~��`%+����3��mY<���տ�<�����F`��x�����UM�T)�i�hJ���AR�k���������WU��N>� �?]�S��^g�Sa�=���n�O6��C���,��3>f|;|��?�7��pyX�(+���������+f�*k~tv���CZ�G�	\�
e)7TuE�aq��l��;�P�˟���732�4]8~h��9qV�YC���u�`g�}v\�����S���AQ�p�W�jz1�O��G��7Z?���_U�At�u��hq�Ũ��ʆ*�Z��E�6b���-	*��F�K��L���c���S=��Y۾������ɪ8㡗S��+Z�W{�4$X��d*���E���Zm���-���r3�n{���K˃��/B���Jg�7Dl@�!�Mo;T��"�g�B�K�jǹ�T����Ik�]6��#������W/~�777\�����>�K)��J7�6Y�=�L�X*G;�;;��X�!��9�<�+�-�u�x����\ʰ���祚s�$��cV�f�8#�AT@W���ZFCUSh�j.�S#$5�)�b�KO�F[��-	�5�'zVR��`�U��+�q����խ�D��Μ7/$]������r��C�b���%p"L:��|�v�_v�Pcbj|P�
���n)�5Jj9����{�����k#�����?���|�o�"��z8m�u
�+%���y��k*����[��a�u��&�`��ϚDE��Y��#��Lיah�lq�̈́�so�ԛRfq��iBAu�ns#��jSiҜ����,��3�j��9�����ss���ұ77�Y�1IM�n���ګߵ;Ҋ�Kwև
L��$6��,x0����Bѝ����K���J�W�n�|���o��[��)���F]3� �}�o��c��]�)�ZcO9X��h�u��1����
�@ur�^s��~4�a��&��YU�i�֊Dv����5w���\�W����4�T%�4�R�s�UEgX��lzԇ��O�/Y��Q�@�s��[��rH�gb{g��I���}|��
�}�-�}���j���(�`>�G���ƃ�P|}{��$U��F��%kQ�����klhF���=�h��"D;�Y4~Y!ns�a��?���wD���&��p<S�$P��;�MUH��z��T��`��/ް��AbOB�?݇t�+� ����,�Jz�wt��u�ŷ�Y|��:�_��+�4�O�������o	+�3�sj�k�R�d�c�)�w�ᜡ�޽����� �G��.*�&#��f�Ki�P,�sa���R�����#�%x���(���&[ ez�R?�Q�j��O=�>�f�n�G���|��z��J���q[e$�����~㼿�嶴\Ĭ/Gy��.<�!��
��&`�y7;m��-��l�B�9(*�G��,�nL�ڧb���^^
�¢Dk0��LS�o�TSo�̍��D�PX���rQ_��O��^�u���]���t��$ `*��40w�B�ːy�Q�/� ����?�[��gQ��OS����nKk8mA��Z}I�ZJ^�L����t�Z��}k�X��_���p}U�U\��g�梅���L��	`d���J����p����cQ=�d�a��s����zS�2c0��Hj�=��Ii�*�=Z�!iX>��������*�S��.��3��+���qL�J
�!ְ�h�v%@@��B�[�����$�Lt;��4�ٞ�(9�N�)�$�R59�����4�p��Y�|\��3����T�8͕��t�{�^�}��jy�V�4�P-���2��R�ι���X��e�e����(��D��H��m���/�	�_e�ZU֓�!X��o
�\KN9�6!̝�
�;|h�%�����K#��	ߌʺ���ٛ�W"���(K~�؝@�o�Y+ƶs����}Mw�L U�`
���jh�d��wV\^��v��6�m��@�Y��aJ��qњ�-Q�~[��gv���zB�ɧ��Q�RI�qQ�}�K������2�}	R(�l�B�fpg.�*���EB�����᎔�ZY�K�vN�Y�
��$n��7Z)�v.�-�Ja��� ���p��ĂX�ni�/��J�b���|����J�����ۧ�9������R�h-d9]���G��F�u4j��>zA�DѠW+| �cڮ�:��LSP���h�Ǽ������I=�k�ޟ�>sߨ-*���ΰʯ !՟��(H��,P���4p6�}-��}D��`��I�Q�cC�!t��M�J���2rfE�`����pt?U'�Y�=�/B�w
-�ƔTi0�!�c���;{�RV~�RHT�ń&���t�/+ŷ~ ��|�t�����z��J蔽 {�V����v�%���#G��a2��өГ����`C��Q�HBs��om��_����=�뷙L�1��9�;�W�� ~�5<*%��t%cN\`Hǂs��4�HDr��+�-akU0U�M�(z�nR��⬋vvA�䣐��M���ϫ[�w='�(��CCB�g�</�¹�u��uFnt��Q���fOh���Q�� �P����N��8�����ێ���/4t�r9�0�Rk���};bk{u��M?��	�AQ���!i��Dbl�g�� �:���x����^�B<6��7�o�<��� �=1-VT��\8Qm=kw4`-�t��rU�s�Q����x���N�)s�~�`�KB�N�t[Й�b���MlR�S�=3���Jb�=����Z��r��(�b9t�]Y�� ����0,�)���33��&��f�d��S����\Clwo{ԇ�(0��HX�����Y����3|�S�s#P�R�,�!��Tע��#����X955���1,L��9+Y��&8����/�iw���	1���*����O���d?�6dwק�o��]ȇ���(�9��k��ҳ̓���P1��gy��<8<����6����Ű$#�'q�sSyRň"�ݙi��o�_
3��x�M�\����W�;�5.���CFb�;4:�E�s�W�W�{�b�׮7����K�3�������7�,���u��G����)��y�3᷹�;ҙ��BP��n��=�  ����Ļ�Ģ��*+%�`�V�iu�,�s�^4s��e����.���Y�lK���!�W"����O��_j!9�㧘���K����N�L�v�q7�f&�',I���)����{/v��j�H���ϲ<`�.;�F|�M6�L�.�sO)xT���Mdx�4z�V���-� @
 z��QF�y�'6�Ik��W�9�3�ǂ��z&R�C��o(E
�Ύ)ʧ����>
z�<�e���^-	�}�,;*@~&ۮ���5���t׃_jp>���zߣ�7���3e�%&�:��,�k|/�a>�m:? y�)�����ʌ �Z�X�S+�i�����#��2@(>����Oa�v)s)�.��)����v�tfM7�c�vH�pp_�B�u�V�w�����V��~?WVT7�s!��P�8�b��Q�� �3���a��#v>&�,��(P?�;�q���vxY���7�m�:�eRP�K�����c^?Hzf#��7|R�9N-vE�����~��X���[�y��N�'��r~"����ѽh�����(�T�i]����r��ǅQ ���U@/I!|��T�ڽ�뫀Yr~C}��~$2Mz��-�֫��L��Q�R���V�E�r�'�
Ob �������4�%�I�g�X�x�W�7'�D���p���Mx����SJA�.a�����L\�w��T{��G���DҺl?������_jᓯ�����JTPqf��|�߄c��O\�ޠ�S�]bK�c1+ܸ:�V>���
]���CI�O�U7A� o9�:	p�X����̈́S�>�k��%��D��{P�G��쟻�*�����3�0^j���ǃ���銟�]	����tI!��4�901�ˢnӠs�cC���8�βL�BW�'�s74�Q�f|S������#���E�;�m>���[��/�e
m�i��T��� ����{�|��RX"y�Tp��82�t͇�/�Rq��>Pܔ$�.Z�q䳧oS�b�A��/v����:����Ъz����P�=1nj��o���-&�>PRW��s1�8s�o���6�C/��	a�~tX�l:ϥ+���@Yk�yv�'���HB��[^é�ogy����U�T���
�2N\��ű?�j��2�x�<��RzBdU�O��nb��Hg�]3���n��M?�z�I�|��'�n��!E�_�;�
H��T⌞��z�O%�E��̘q^�����Ė��1��\��+u����PPd��x�_k� ~��q���4�fds��d�d�A�QB�W8�8��Z���J�N�#J0.^�{�];�l�])� `�kx�"�^P�3�#T���q''�` ��yH�6��Z2_�* >v��ږ�DST�\�5N۰6��p�����M·
��!��|n��+�2��W�tEY��=#��%��_=��L��.��do�6�3%:<�r:�6�y�i����c����ali
e���z��E�=����K��H\��aZ>HỬY�v����8��J����%��w�=��YN<�q�$б1���L�gp�,�^Ω�[_������X�`����q��Fd�ӉO�-�Ѭ������3_���`&/_��ȝ����C޴qB��h.Z5pm�K���&���;�	��V�α�_�z��_�ru�LT�S�S[bߍA�L_)|$-�-K��&��������Ns�N��oV*\�m��ʼDe��ӝ�&����?�7΁�+��ղ�H�0>�
_��y�8̫�
x����{q��`\�_���VJb/�z��ں|�%�"��7b���C"�p�$��c�G<W�M��^IJ�sڏ,��e�cX V�1���q4�E�p| ���p�A&��|�s_+8�� V5�TJ�y����`��y��l��_�I@����s<Qr�qO�uX�tt�w�G#���
e�檵�f�*ހy�ޣ�*z��v��P��c���3|h����_����}���{ˏ}�9s�ƚ����n�̿ӟ�*�al�%^��oPU䑇|��L78ҔX7�_�d�py9+$�{��r��,Lz�I[����y�^G����$�9~��K��wj��i��$p�o��;H��+�nՀͽk&0�<���]v�}����7��g+�Ӿ]�Pa���(>a�F�h��p����فJ�����Ҏ�[�H�^���iR�bY��+7�cS�����y`e��aS�c��g�9��pK'Rt�Ɗ8��W1:I�2�0��Q��J�I��ʠe�y?'�W�ٌ�@$�ӄc���p�H��M��d��h������c�ۢ�rW�p�
�(�b7��!���:�&BѐK�y�n�^D�Gj���b֏��E�)�A��Sq��]B3�Y���b��r4���ĵH�H4?ˋX��Q���4�b��s�4f{Q�n�I�a�"�춿�w,=,��X�5��ѡ t�kdr�X�\���)�:�����"�2L��R��p�����u+{��	��>P��X�֝w��<���
.�6VH�V$�����Ν +����^��:�fW&�C?I]��n�Em�@&Ւ�E��_`����F�v��-w.�y�[�Q��w����ؽ�3�V�&��2�o�2�y�ZS�Fj
�5g%��m�����Ł�5�wl�C�MÎ��;013������R,�.�幫���J��{x�H|�N���^Iic�Ptɋ�i'�3?�Z��W��=��Ѻryq�r�i�w�Ǟd`kg��-R����	�����e�����3OcQ@�'Q��[x�5���[@�-ܺ秫�sW��hҍ\]6*��2�~w6Q��aJ��$X�qd3�A�1��RQ\4䆢��ݤm���%���*���0y��T�N�!������8V��n���Ii�D�>Ӡ��#��V*n��X����B�VT���sL�����yIr磃R���nf�� �fj��!�w�����B�!�Dֹ�
AB�0��K��؊��j���H��sC��l%�Õ�IL�3؍�Ő�|k2'j�����ҧ(�I�}a�����n��|Ŵ�d�����EL�����G�m��^~�m�Lv*R�2�\\Y��m�?��q�#A���;�k:E# ���/��=��/�������x��0�s�^���1x�/���vE$��ʀ�����i.��y����wI\]�o�� \�1=��^����8zH��y�p�Z�,D�!��`�J��>}s���*�o&ؓ��0ױ/�_���A�J�5��" ��ʌcoWj̣s�E�� ��ҹq#gj�,ڗ�M�j(�������e̸��_Tt������m��	���;�Z�w��0��)j����DW3Ie��ث��h7�����G2���Tr�s"�m�W���Xq��<�|_�B��/�r�￝ʛ��R_�f��[�}��z�D.Hfs:���̥�+�Ck�+��R��y!��b�5О���TPjhy���𶑯�2��.�/�3&�h�5���(&�=ۂ���ԙ�}B�9���zJ
*B ƶ�"*kƶ
<����~b���MڗFN�іAz'�OA�,�@I�<ጞ�ԎK��y�ΛT�A��#�is�\���"�E>;w�Nw�亡+�S���u6���P����P2�K\�g.8㩸ʙ��b�}s>< �O,��k5A\�%�*j;:�h��pf��C�s� V��:v]'Ή��l�@�
��C�����������P�����/�U�Յ�yX��e�YIw_e�� FFrS/F]�)<��`�;ѐ�S�f�[,MCce����nU6#,�Bj�~�]þ��qOG�z11,kӆJb��&p�~8�����H!�Ue����趸�˘��dqY��i�"_+��rx&M���e�w����B*��'��PWB�nQ?4=�y��1�w �,P���R�b��$�o^�2�_�V��s�����V ���y�eC�1"C��K��I��\�u�Z"��ޏ�; ��;�Y�q�m�x��×�ns4�L������锛�������s=�%qA�)bV����D`������dg'p��*�J�QZV�:^�Z��~h��.���
Q�i�/F/
3����[��`�#�~Uc��pu]�l�;y�
'�3���u��h�h{w��w����._�S��Ju�'�A�[������f��-5��Ib����	��,.'T��b��54Љ�O�f��rs��Os�o(��Qm����
e������Z�s�Q\{Sd�(	����Q���-VoE�P0�i�-�M^g[��� �l/ג�ȡ�E��G�R
SL\?5�#>��a���Hx<y6�wk���u��Շ/�z�������53�%�s͹��*a qn��F���G�<�x�a�9���D���f���m�����3�p��l2MkAS�|_�h�ǎR������Ј���i-H��0�'���=�9�q�&h��!�� ��Bd����cc��~Sd!��m�5U����`:2��-�� �5��i�S讔aņli�@}h��^x�,�1!� θ���˚Lb�L٦��T݀\���,)�h��!�A��	�h�����-A�����" s���d��1��QQ\3𰘘��L	����S��-�M���DYݖ��KGO���3�sW�]((?<{WG���L�쩒(䮨!Z5av�b[e%(h]�+�&0G	X1{�h����p�O�6~3�Y��h�T���狺��()��$����y���܇�A&g�k�1�q�j��vҧ�B��Lm�����Z��S۠�&�i��Hf��kĺ(KY���uQ�0��y�+� k����ۊ�� .�L��S`�J��ޏ�jx�n:�LA�����2q"	�Y��/ȅ>��hʧ`Sy[�&V7@�}�\_D+:��lK΀��Z[#�)}�J�k�#���7n{"��j�P��̯�~�=��&����{�YM��:���c3�'��"�Qt]lo_y�K|�8כ�[��WrP�xٔ��!�}���+L7��^�{#�3KX�%(�s�V�"�Ɇ.&@.�ѕ���%�)3&������:�h820m�g�Ny�4Kt�%Ûd�i���ˤ��U$�]֑�r&�:�"��9}��ȗ=�K��//70)��f�U�� %>m���yF�dP�j%����{&с_h��XP}�R���9En��2�wX��D��ك�o�j��s@�tL�@����߰L"qТ�}Ĉ����Il��_�NO�Ĭ�>;����
��j ,xKY	��-����_�cXac<LK9���| ���A�y8�i�'Гc�bzr�G0_�YkY��N0Q����	n�	삀��Ϟ���$2�oCN���b��9��*'f��!qY�����">-�"�w#cy��$w�p�J����_�=��~��Ų�Ʀםi�f�B���J�������hh�i��~��d�Gr��R:��1 Nӊ��)�Y�u�L����JWdϯ���Wn��j���	�b���.Q�	��G!�ӷ�{ �����s���V8��h�l�(�(��@ςԛQ�z��Z�I_v�ZU�\2<յ�5����<�QeS��y�d@;�&��xeD��o�t
�����?G����F@�������G��z��.�����EV��;&Nj�.��]�s���P��\0��s 6��-�����=Y՘��D�,��t���:YzEh������=;A���fJ8�7R���=�c��\���7�ߪ�Z��$Æ���2�����7}/�  ���{�`�>��HD����h����~M�k�����U�67�A��sd��R}e���3\-�I���@�[�)�fb�CĆ��=R���/��̄�vwA��4:A,�q!����, �Re�2���M_	����2�\jk�ނ�n�����?�iT��������2'uMd�C��LT����@�pF1X���Ͱ�ߦaEQ�#��{����Ӆ�R@8���u�Tu��݄t
i��� T��Nfd��#;'���+�sd��>�:3\N���9OE��/����*~��9�N��R:��4�z�%�G&Cѐ��ph�Ȗ{�/�Z,�M$����g�����9zZ]9�.Ju�72��#W�w���׬����P^~���(t�g�"�p*�������?l$Ӳ��i9b����)`j��Kѳ��4}��~���w�)n��w�������S�����2.	w�V
D�� ��֣��|�W�D�D�[����/A
��R�r�pyJ���]2N�4�u@���$&@�����{[e^&���_�p'M(�VkI8�#n~�#	�W��MV@k�ϋ@������J�1y�ah}F_����)po���
�s�^d�T}�!� #��1�il�� ��_	��-4��Gω)�q�Ykfl��j���D�q�?�����\����v�Z�I&D���;����=����xB;��*8tЅOƑ��>��ۅ4�*80U����M�#�u��� �ҿ�W۞�)��`����'�p��a��\ǥ��G��PH�����'�������#���QI|�k��֌p
R���5��x\��M�N�\j��u!������H����-��w'0�d/��n���w�؞��Hsn��v�7�_��aP�����p�{��4S"�9{ ;�t*���m�1S�Qz�j��t��89��뭃���C>H �$�F��c���=��uWG(`�ȉ���pC.M��	J�IG�_���[w��������J%�F(BT�ܪ=�쥡�~�-p��+�ߞF@X�*J�o�O���7�d0��>��a<N�ްѴ�O�,;�z�{<��T�Y���}n��4�39���T�Xy�Ao�
d���W.��CL�ϰKc��S�k�	�:,�� �0��Z� }�p�-����n3����w���x�d�4���20=���A3�p,0��̃�ދ�:ҍNo��Q����3�"�_�V���P�1R&�g��%�B�p��#�a�!��!��0H�čd
`h�u����7��LHc
O�aAR��4�A���îa��=�D��nr�,���qW
��������=r�:��f ��vrP�V����o:0s���]C�@�S�Y����,ܕ��:����4^��q����K=�L6�i_}��g�<��8��>yB���P��ﾪm��l�$�rM��f�b<.��9�޻���E����Yl��
~$�{�h��i_���L�1Vw�3��^�kN
��In>f�\�\��څ@���2�ퟍ��������|�/L�?x�j�ߝ��RM?HOߍ�K1���!r��n
��ϪW���%}|G��R�F���Se�#hY��_��d��JR:T��w��'A�5�S�;*U��q�x�I|���-�C��0��I�R���������ђ�����S�
2�bC.��٦Ma��B=�;'�4�4����4-��xt�^�������WԤρ�w�����1o?�Ek������Tʲ�{T��MYq�12yM3o/N�wD΢�"���	ǝ![�X[	�*%G�"�bR�Q�J
�#��H����4��"C��"*�&;g`���S�MsUY7�nL�*�]�m/�?����l!�����Whp���k�� ���-*R�����?G��5'%��݃�E�J�U4�
0S�-��H���w�������|����v�K�b
zJ
�������Y��8ӱG���l{XhF�^(� B�e>�]��K�חƂ|M��������-Y��]x�?���kU%�,yl2ew�:�WYl�{y&��k3�����!�	�hN-�TQ'��z�|�[��n�s��l�=d����kO�d����[(��m��	�ң�tD���m���ڷ�5�
�92�R�ˎ��y<��V,d������6w>�^
�>����y2�$C��$��������=��jw8��>�{>.ƹp��&��V�u�>c2�:5�G�Q#�h�q�x<�T���M�]�@�!��P!7:�� )
iBE����+��i%\�u3�0x�e%Ȅ�X+�-��]��~��s/=�X���W�%���V�A�έ�p����;��\Q/����J��Ցt�m��о)z�Ey����Q.�x�s,osD������h+"�+�a��K��8s�7�<D��s�m!�/���|����(=9)��,f��3/����8ܷX�*1�S�/��65�w���%�zvH#�0�H|v�,�u��@$�S�ː�C��ɥ�����	h�D���Pv�4�+ʧ~J��{�v���Z�[:cQ|�D�ܒO^��(_ ��$�D��d�)���$Ѽf󒼫�eU��N���ǘo��6I��K戩�M�<�W��¡��Y4�uyV��zp����G�^Y|�ԍ�Y������,cSK�M����[�� ��ߵ� ��J�z�Zu���V��:�];^� ��y���^�eS%�V1V��l�P�PZ�fL_T���GJ�b�q��\@c�n��1o(�
�0 �r��!X8�����<��<��%ZsT*F�`�0���+/��\0�Ր��"=;�S��hKgEX�7�9�pIW�~���ϹBܮ�ے��S��h$-��8��rޔ�'�A@b�~<�u��. ��F@F��vx���%�F1Y��PFG���q�l7|�*u1��S V��z�L<��<Y�ԶRp`a�[GiqC!/y=fJ|�c���첛=�o�i`�����G�����V��p������%���A�r�ެ2�n�xpV�d�&���z���(�e�5����j�����8P�jOt5	�8G���`���EBj�ˡf��+�cx�+*��	�H' �B���5�Bv�Z��[��+��c��i���n�����(E\��`#��r��9�2��¨�6�1LE'0���������Yb�����r�t8����Ֆ���nj>�'��C�TP�����A���'b�
�<c�|K�
D�B\B�G�5�Ʊ�|K�n�aUg���K� q����U�It��(S��O���l�|���ށ������L6G�}�V&܀	�~
ZZYF�41�$�#�h�n.�������\0��y!�(�g��7#JU�xw����o�t��e7�]I&�>���BUID'���R�uEJ7Z���<�t�6�q���%R37r2��L<u�M�)�p�#Y���9����m�@N`�W"�����C��@��^^������^?�A�g�F���Բ�J<�W�f�vHa�ͻT�o}�-#v��w��Z�����\�r�1(r.���N�6�����e)�k��yF%_�&1�=	���I�3����ϊ��Q_�g�>�1_*Tk`�Qf�0B|�p���BFTR�JJ��q8��c���=�5��c�=�ko�����`�ҿ��?���߱�M�:Ҭ8���P�I�+��GI�Oc�f]�X�k���]
=x��P3O�;�3碘3z�z��V���1��Cd��@�ʗ������� K�dͤ@�\sffeO��Ĳ��jj8v��./�p�0ς�_����N&.:��r9��or�F�͑A �z��F�yjb��H<���P��٣c�oп@�Bf!yf^��*>���O� ݄�r�t�f����A@F[�l\��L�z��}E�?
�=z��<1��X�(�!��j@��O��I��5������鎣�@ Dˢ����j�$~g�<��.P��J�-m:���gv����L�;��fJ��V-��N#��u�)�(�2�(�kX�Î?I]�?Ke��G�+��]�`���{�H�7j��:���wx�X�E�/�f��i��E;�(��w4H[Z���.5�uJ�V�3�X��jê������J�����Y��Cs��ʜ)'vs��Z�~wvH�#f*��~�b΅�D�iO� ��ҁeȰ�4�K�P��y��Q����ii@���98-��ywf����/��9\௼���j�^�����[�;?}���M�Q�^�K��� �����Is`���-��f>m���)Յ�k�J� ��r��Z�����*���ћd[������m��e�k|\�b�!������ƟW�2 r�v��KDiGy0�=G���l΍�J��s�p�ސ ��<�u3f֯�O�>	%���̳\��$�*P�<�׸z�LS���})@�E$I�ھ�'2iteo�uK��wuI>��Ֆ�OPt�e�*Y�+��n�� �ܲ���ks�&�_��(S�-ϨD�du����EE�`k�dʀ^ӂ�a���z+t��4�M�8�$w��;�?�;��Sm�7�.	U1���}����u�;�-yl����T9��R`?���Y�%��{�M������Dui�@�W�2�9+���� ܻP�_䮫S�-���Zg��32ݿ�w�@8,�X��y����ꁮ�*Pr�X#�� k��=�I��
:?�E�ԨOo���0# H�{�u�WK�0-r fؽ|=!"8�١=��q�|�݆J2%c�`����f'Eyk�h	`ZļT���R��n�>�H�I�g��JU	J��g�ߔL�^��n���zw���j+jn�ep���O���dtsq��ɪvYR>�:�j�ߥx�������<�.�x����齃���yZ|c�tuJ�F�f�`�_��W��A��TW���m�K�C_���NݟhK��d;S�I26����#��@Xhu��Ʃ-���N�
�fy�4J���{��/��i��^��Rl���]�Ɯ9=��Vh�e;�}N�r�Z$uϯn�9�a㧼@�KHG��#�28�b�?��E@{ܙD��/h����H*�z��7F��`���~M�F4���mX�S
��
�p�'�!EJ�a��d�:��HO�[_�s0�tfnV�����[�C�������~-
��P)����Ғ�˦�2��VT:��h�~҇���.���T _�3��6�[	����U�&;���-a�ҭ���D�Nu4y��RYw
t���e��`ˣ�B@��|�����P܊Xe��5�2��;;g�D���a��s,-4i�B�
f� ����5��Dm�c��o ��C��6e��!i�Y�e��Y(���]�~N�cs~׎��q��z�F��$@�Y���ݯ�U���ٶ����y�Ft��������H��(al�=�$~��A!E�x�"]IX�°YRE�mV�<L֒h�H�t��j7B3����QA帯�Z��3 �I��ڡ�p	b��&D=<���؍2��������b �UOv\�	4�����{�(�������Z*��rw�l$5���al��h��BC��H*�t�mK�D��*�;�~a��}�&"r�% G5����DYU�l�_\ə?��L%�*���|��EY�`o�[��پ&ؤ�*�Q���θigM�(u���;����D���w"4�ϥ�����fㆺ������?�\�X�ex������@u�\�Ȓ���\�b��S�Ä:��L��q��3Vm"U�K
-yu��%�����"He+��*aHH�����:����g 2�f6t����hB;����.�l���ga���O)�3��+��d��i����x��$WQ�nOL˩��0�A��[��j1ގrI����}�.��?�����7[������ϛ8!(/�Ɣ|ˋ�rbY�%�1����]�d��NC띬o��>y�s���N4X����k��;�v,�4���%��(,�G�,�Z�/G2c'�k;�OWN�p}�5C�gY4q��nX�q�l{��o��&؄h�������%Ɨi��w8���]�:�]�?�Z��\��no��E�����E�v�xf�:���t����$��M�5Y��eG<�Z�N�2{��7.H��|c�����5m��UM���H{4}���_�u�J�f�h;o�b�&[!$�����%��0�#ܙG�q��(O�D|�=��k�o�B����B]u��v5�|�[�},�J��!�~���g�o���Tn�����6xM�{AhS��3<[���rc����~��M�����Yb)/+��(7|9H����n��%�L���q��9��bR�s�s���Џ�2Y��Ln�h�(vK�����l�&�B}�}�ip���UZ8Hlt�g�K�e�}�zM���qLAq>�?`V�����2�W��T�3�x��	�9����.�ӡ�	L	��qQ��eu/�th^�[�j�m�ͯ�����w.N���t�+���@�:m���	kY� C���&�3���c9K����: ��(YԶ����Ш�@;F��!L�4�Ml̴������c�u[��,h�wq�hCy &���~4\���g���f�x�����/'��h��.9�u4o�%M;P���3~~?i���&�-c��8�3]w�
(��6pt���/��)s/���K"���~Lq�#B�Z)$`�0Ѱ&�%m��|\1(Fj&-�[��p���4���2L©�wQ��Uo1�a���`@�� �!
��х��^���B���X�Z�CR�-�t�Y��=Ks�o�����<'�W��s�|��AOZ��g�/�	7��-}km5�GK@�ڑW�b��XE���~���ˣ����U!�~��z�.0�6DFLɸ�� >ݞ������<h�A�������T��1�R.h�(���;�P=��m��:��Ն�l#u;а1҈W-����i���#q*�X�c����O���"d1���	q5Gt���F3��K���ꟽ,�$�42�����"�Ӿ웛�������|h[��u�>�;LD� �j䡕�'=�
�I���b�z~a�c��$Ҩ1��U�m� ���/µ�&�qhd���ٴ�2��&���:���[�uyS�D�(���`���#.�\� ցK�m��F��a�;/׸r������i*����=`ғ̰�/��b����u@�a�1����w�_�F)PY
����KM��|���g�+�A���+�;?����M�Ml�HJ& @�d�}�Q6R
�ӎeP�#Q��g%��N,aI��2"�x���{�PQN~�|מa�\�N����%V>̕��%
E�&R�ƪ�!����WR�����0ߣ��%�x(M.j�XVy��&Q1Y���q{)���!c�d�WZ�
3�&\k����:yG\��Ci�9���Dr{!|e��u�f��c9`&P�x�\����C�D������5f�q�e�8�r`�ۦ�+�]�n�S����d�ɬ^+�JQ���cرt��3�"��! W�D
�.p����p��'rS_,�R��	�W����DB+�)�U�@f�ۖ}��HJ�`������*A)���_��� Ewu�A$�:�Bx*O㋌[�C���?4c�=s"7�|�/�.��?��J��}Ƹ���9A�̈́��v�B=�&���H^�����"��̜ؖ�Atm%\�"R��H'�TP�J:��	=h�p����Y��(~]���
,& a�����Bz�c[7���V���El� o�ֵ,���h83,8l��Ͽ� D�tll��Z������b�ϒ�}�i�"�u�����N�L:h��aD>4�����b� �N�b�;d@M��{���+� �]�8�6)�Q1հѩB)���y��a��7��|��#��n&g����ɻ6T�������~�Ϣ|�À��r~i}����#b��Gx��}$	]#�����wjQ$gk��u���A
�G���,�PE��8����M���#���~n���Hx�Ex�:̗���-]��S9�a������rOD��D�W�[ 6@F���88�b ��C�X!���i�d�	c]�tأ5�p�y�_������JN&ސ����4�nd�����������Z_����c]C�;����*�K�zr��l^ؽ���f�7hf��c��;y{�&���u�lͱ��p�� !m2&F�u�L$\���BN�E�E�b)(����[vn!���gL"�/��mM�?�,��j��� ���x�;�I�%EmJ���L����4�b
���ҌH-�Ѥ��&�&�%g]��K@�9�|I�璉x�s�2k ���S����b��0����A�r/P�&���B,⦐[$^�o���3w��o7�������T�$kz�t��O
�+��7w#���˯E��V��b��ϺoaV�D�0��ƔS�.���e���5��.�I"(�_�OlpA$~��݊\���D�\���6]��}���}��0?eWS����;���8���$�iͅq�ѝ���Ȫn�&�6�W ���B�|�fd��X�q�7�xB~E��.^��/��-_4����QV^�Ϡ�	%XU B�(��/�z�nO7p� gX��Z�]smA�jy�/���]��[��Z��N5�i�-��U�&���f��),�e�(�Z�Fk � �&�}Md�5�Ude�'o�7�})w�^#�Wj�Ւ�_`R���Za�nz���V���g��A'x�)��%�j
J���-���M0ףqjN�T�L�KmXE� 딪�����2p+��k�n~^��j�p�<�'z�w�����x�c7�����햻[=��v�/�Y�a)�n��&ۇ���0��;)i謗kw�h>�9f�}�Ϳ�e� ������d�t�gU�� ��t�Ѹn��E"�>�e龽�B�4g�rf�'��U&�k�_�� �lG�Gx��q��@յ�p��F�+�)�j���1aw�oF�g��Ơ��GCQ�"��1o/A��s���a��@���%[�9�u��'C��2�WE������UG��~�J��Q5l�}���J�N׽��Y����ńP^�.B��Q���� Au,AE��!��5��&���ր#��"�T)�yIF���TH��L���z���9�����*�>!R��wi=�}��xE�e�V���H� ��I�E�Ǡ�Ͻ��zL]:$��}E\nS��[��EL�va��C2��ғ�ROwT��vk�>���X^�9�j�jq-�|�\�n��-�w[K t)1��nIO,��(O�R��}%�8��=�lYV�?�7�q�&a�-9,�ɬ1���2`�,���&�n�;�r�Z�n>��95�꾐��y�H'ډyد�����jjE逦��+��Y�W�d �~x8P�NB�<�it���<�i�8@�6��?A����ϫh_Ky�o5�HvM�����-ԛo���Ӷi�]��^pn�hj�I7�����Pr����L?}�g�C���v�+'�q�Z������OV�j{�Y��}�5����0����^�.b�D_��[�\)�X��2b�S�5�cP7F){����BS�6U���6S0K����p����p.Ρ�v/1o����E�̘Iq��m�J��`SE��D��*�Tv�&٦ ��i��b{�T���<?�� �ʽ<�K�%�,�'���^o
�y7a��ϔ��8�Q>߳;�?3�<Yⱳs2�C�Æ<��1$R�s9�l{�ԮC��g���?V`a�4E|Y�3Ξ��r�W.z
A[����2V��K�CH��&��%��S¼��6���,���ū|�@`��M���Pȷv����r�����X�:/t��A9�����{�kr��=o�D[�*��"*ı��&�K-x�=�[�F�f�(��H..��aD�!j	�1���n�V_u@��Hn;Go؊��`�v[��ϵ<a��)�g�'Hˉ�`T�z'(�9Z�;�IdH�+�T���f��y\�pK�AI�^��K�΄lz�g)�����
T�_�����l`b�>)���ԥh�iħs`.)�}� W���7�Խ�u�b0�J �C��f�^k�=ѹ
�#�=�!��͵{ǚ�"�.<_`VT0�%�:恿aY�p\D55��J���)y�-K83�@����VVۡ���&�	j}�p~6ҹUotJުG����x���.��P�"(�!`��!�_���eID�ݗ}�Ҝ���M��q8'/�MTR�Α]�$���W<-*!�N��ȸ�#�����Y0r��_c�?h���n�#_~)�@�>`6�<	6>X�?�iMp����T b������)�s�|]�8^�$g��^,j�0I��� �B��%nEl� ��,����Q2����"�9JQW����$6G�Mb���T�4�i�zg��p$ʋ���гk���F�j7���M���[�� r�(��=5�ج��Y��}��C�L�>Td��z�a�$_���q�/r�F�d���\`�ugO�k�yW%ዡ�xPNگ��fr���P�u��{���#j-Fo�ⲛ�G�iV�	o�C���Pb�M�# t�V��ř���(�c����'W/o^l�r~�%�/{��h���w�yش�|0@�;�g�@"	/�xXp&$fE'g�^FBTĐ )-�
i�ϥ�����^{���b+z��7B|�
���}T�F�ֳ����q��n��+j �F��}����Lev���F�W`��E���.�n��|�42;C�D�-���%�� ���Ĵ����֓g������u}�� ��%9'F�/Q�ɭa��<4c��=�s�$��0�.Z79�^���\�;��d����(XS}�\�q�.JϦB��e��b�lE�z�u�Q_ۢdmB��>�!�cI�4S]NP��F�y��
Η'6�X��J�5��jG�x���bZ��1�Mj܁i�D�Da3޾���O�����/�q���@1D4�7����m#�펮�����8T����{�LG�`�����Lm� Jި0A&��^��[�0V.(�@}��9q���Lܦyx�E!0��JP��n*Yd
`�ICR�_��X�-oI�n4�f���0�Vp<Yd�FPI����O�vNv�/Cؐ�� �>��c�s�kiY�-�IB7_�L��rNX�X<�4hH��pЪ�!�õ���:{��9��P)ྡྷ�m��c�/����9��.r:?����۽k�eJ1�kX�;]	�S7*7��6�]����k�Xi��qړB\�g�Nomc�㍤!��|�l��W���%(�X_��*gG.���W"�Щ=��e�m�S��
�#{ά)|����C �n���G���sILe)~:�Q�<"e�(]Ѹ���u���ʤQ��7n(G+Ԃn�s����eI��<_������E<\��E�LE��e�K>�.��۫��Q�4?"��2Cg���h��J^VVWf)YmzXt-$y�2	�_ �:��	62�ss8\2�w�O��fT��w�葙+�
 Q��R��vna���i������2@��U6�0j���2���P��^OV(�.��v��>;E!�X�d~f��v�?����G���z3����x������hjy�9��^�$|�]ָ����3Z�s�q�֦}�d�߻2*�303�X܃�(ЙX�ó����by���k�'R^,?�%�k�D��N@�C+��Rs�٨�P`��q��h%����?��`|�d�[6�v�������d�J���P�ԩ<*X����*ȿ�~1$Kl4 �\��&����? G! XA.��pZ��	9���/W�I�c2[(ه_�`�%j%H	m�N�T�:�K��й�S��|�%VԞ���p6����L��7�=7]��	Jz
�L��w�ԍֻFa&���_��^]������wo��̵�1���l�o��U��3��m��|>��(����X&�a�π�u�(�X�M3���Bٱ�ǋ���t~��&�����Q]�C��壊�����m�A��)ľ�i����t\��	L��_k���#��8wh�����Z&V�ye���j9�}���x:Y�&�� fn���*�u$���\4�Y	��`�V���ļ�ƭQ��;�"���f���>��eU���{�E�ԙ)l��A\oԋ X�̽Ln����T/��ͫ��gK�m�u��ڭ���������j����"w3*L�tq����Dٷ���;D"�7K�]`�B���<���p���̑�A���B֋o�8��8��׾���)���9��vz,�Fw��<0FlP�UEUAf�oFkۗ�#�I�￻��n�$�<_��Xӽ����������m�L����]+@�0*(�8@�a9���"�����x殌t%���*�0�t��`�\69E�f8���C�țDi$;6�{P�Ú�IU���c~Ú������cx��$*���҄G��}�ߓ7r���牶4E���뷨��2����#���[{�P�6=�V�����r2�M���� ?��et�~�Э������k[𵷭�Be��*T�fS��N����s��Z��>��L��X ny�nǧ����=��>�
�w�}��o�X���Y�7yr��Ƌǣ/�i���Y�ƻ�k��LW&S�ٌ��_�(]�"�C���:��|���\�X4G�/|X#�N���k���!�ۏC��\��U�N!m�,w,;�l���0 7��ۉ��G1|�]�K������s��5�g�܂��dp��ꄸ,(�֪�=1����]�,#~��
��)�]�Oq~>�2�h�$Ȳ�yCV�.��B���uy�z��;�d:Ϣ�\�[�����B�C�@�A�J\@No����tp�Q�:���
D�6�����~����C��b�:>ڈ.6>t�\��B$��"z
�,`��'���(�#���7�����n�p�.�3܍����e��պ���L���ʤ�ߙ�R*�W��~��۱'Lއjed����<��_!`!��x�Y�S<3¡x�7$F�Y�_q^��f�˞�7���h�����%��K�� (dWܹ*��\����x0L�y2��j��K�i�m�j'7�?�M���\��|��o��YO����Z"����a�j��`M���ڥ+��o`�'�n�(Z^��1����<[S5w5:}d�SE��|6�^ϝ7��1Pp>�2)��-�mA����{��*^w�[*~ŉ���0K�
�8\c�I X�`�p���`�-�"����#eo�9�v�-|o�)��$]���1��1`Q����s�X"��+e�E�G]�ik9^=c��g�+|(^�S�OF���^�7��U���M3����_s� �d�HTۼ��h�ѧ'Nɘ̌%.�q"��
�����0�H��g�W�y�˅%��1n���߭��*�5w��ra�b�չ��\βy��DB�D��y�Ƈ��՛���ci%y��ص��ϡ��M�d[nQ���*ư�����p� ���s�Ҹ'�Ƚ�T,��Ak��T�I��/\��8oV'z.�K���j�p�w���Vb�ѳ���΀f����z��jY�A>LH1������m` �7)$��6wW�,4��PC���*�f�@���3���-� �$�������?K2E����(%��`�=��N�YfP�T^�� �������[㋳QB횭��7ms�Ǹ���20K����5���jG;Ss�F� ��h��:r�J�.|P� 1�K��Rg�д�T�jw�h2?F���&@�d�35�4?e�e��~����ZG�MR�~���m��O*��l�?�?mq.V�J��������DDӌ�G���
(�/#�d��0���%� !�[2I��Y|Қ�~Z���Lp�5���IR;�o�ڍ�!�QjL�GD x�Q~�oB.e�W*o�U�
@�Տ0���5՟Ʌ���ٽ�]5�\�GjQy�.�Ҳdi�~fZaq-�':� X���\E%q	@����'������HMÙ��Q����������!a�>�T�[���(�~y4c������E�H��HC2 ��>�X�˃5��E1������é��&!�D�^&��<�!@��'�F{�v{��������v��XJ�bC�V�}\�����1r��P��0��z�b�q[.�(�)}u�y�Eu�)�0�/|�|I
A�8�ϖ�9����8�p18�>����V��+���fSX^E�X]�r�����@9T�x�2��ĘO�����P�����2 �R��P��į4��C0j���k�QO	��cP���[N�p,/�ͳ݉+��{�Q\�+�RU 	����]7���LZ��8(������_9���W^���� �G��w[6�*�࿎4��\�x���Q�Cg�YS���B��x>�QaɋV����2w�x��1�0�j$p�}(�0ֽ*��Q�
�f��F�ǚ䔀m��t��W6�] ��� D�Bd�3{�!����<��F>��Ob@z>8=i����T���t%,[t�Y��*T�=m�����+�4;.w�C_3����E�\02"-#֟��?B��d2�Ԁ;X��%�� ^��zg�i:5��U;�d
&zсW:"��ҍ�?g��.wx�֧
w"m�e���vу:�%��D�^W͙�s48�^�
�)��b�mK�b���ޕhoӬ*[�~�$�A@� ��Ø��7��𢯼�!����Yz�ېg�8I�� �E�{9I$����]o K��U3��*�I묍S�L]���%.�E�f\�6���v��ź:[����������c���^��?v�%F�t6��~�\��P�*����LUy�;:\�N
Vt�%;1�|0 2[k޾����\DH�ec_KF��^����Vv
���RsZu�yAb)nn'����ʫ4;��=�^f}�j�Z�W�!�w~�5I��l���^{zؘ9H�����f�I�+k��D�lX��T�S?��Ŝ��[Y|��sc�����<?#����x����p��ד��,����vY�S*�G��A�&JM�Ι���D?q�M�m �0�T��mY=�pg�Z��ل���s[��3͐�G�a��{���_.��>�Q��^Vo��&�&���_nSN��T���2pRp �b|�O����ŧX=�C *�<��:Py��qb���LO��O�^���,���&٣�a����	�Ex�'l�Ҏ���x�VRM�w�S�G{.�&t�����E\^t��i�'���Ձ�K�H��%��Ν���1� H%�rt��`��F� �/sj�X���K�VC��lb���X�U衄�U�Ѭ.)tp�|�q�L2ۍ���|�5.=~��3IK�_?BU*��%E
G�ax�jiQ�y�h�X���eg���0�����38����u@��Ο�$�	������2B�΂��/61 �r�a��"����=qP��Q꠿��H�{�v���i�R��])]���攱R�!�9��-�ewc�����$�b
���%77	Y�ϝ4��F�����q^mH��ٕ1�ˊ�����A@z�������[$VKv#{��YL�6��������R�Z�(�s,��&m�Ep�P��(&�c��e�/휜�JU@�����U��Bv^M��R�Em~=���6��L�˱�0Y��4���L
�A��<?ɫe���E�CQh%{�q]W��j�"��J�/x��c��=|6�x���^��+U)ǝ3��3=`K>D���1�q4	2�b��%���I���S9��tS��r��+���n��핍��ZM���Qb~�Xo�MQ�ޣ��	Tfq��<����=�N�k' �͸� �`��^[q��.0G�|16������J�f�����i)�lD�\�O �5��~�� �D�b_L}�󟮭H��9pݬ��'��W��J�V؏�o�W|�E��,��o��	��Ocun��X����q'�)H�Z3���l1�#<��V=q�bBǓ����Z[�z*����~1�h:�9P���6fJ��w�b��������'��51w��1I� �T�o�.�$'Y�i�j�DV���[�\�^=�RE@����wYA3j�����d�e����))�x�f����o�C"�)-��P �<f ��c,�Kڿ��r2��oO���b	��:�����`�ճ����S��~����z�K��t^f���z���U�J��)8aM�֫&t�rLa6]%�	���Rsо����QI��Y�2�P/�m�*��W�_E�	����9�=	#��-8RP���[d��0�v�.	_�<X�e�^��G$ǆOE���=G�O�t�]��CQ�G�L{�2�٠L���0�^Q��IN3&�mグib�,K�\�ϳ�I���LID�H�~W�խ�r�F��aU�u�/���tp�V�Ր��p+�� ����e�W����.�`,����	�K&Е���Z�u�7�Y��TQ.ڦL�'W֊D./��V�L�����<�����&q���%�1���|��2���F��G߷�W��Wؕ����A����̽��N��-J����������&8��C��n�p��쑳�3�����+������ڒ�BI�!��L�������k.��ǼJL�h�W"B�Zޅ ;JB��%LQ�=?�#/X�뤒��U�ȋ�s��Ï��Z��~-�X�{_w�?��xM���!%̀�(������� ш|�Aw�O�|;el���:
���B���p��C~1o_1��'�n�g�ir�Vn��1]�?k'�st��8���*1�2��M'I`��~�0ŊI,���b��
�l�!O��PT]�tV���
~�E�F����z4�L�L*�op�_X>Wu^�k��lҿ0��{o|�c��W���Iݚ�������HgK�����2��bW_�,�����
Hr���d����=�j�O��.w6u�jnˈ�Bы��%O�dY�� 8:�oۙ�R�\�h��_��=�"�&��el��hV���ol���'�@n���8�nW`Il�+�I����,ݭ>K�bhH$l,�jU�G9=�	�%1oA�d����\�]ം���Ŀ��򀳕��3�h0�C�>�4N��}dq4�������H���t��A�TA�����\9�X�vZ5a���y`��Y���
l��Hqn?Vp01�\�h��e|���.�o���������k����c����M�;7�����f�r,���P�\�`�F7nO����HZa���X���W���$�\�h3j� 1���ܺrؠ��t���g�'`�F�����W\I��4�M؟��yr��*�����b���X����$� �q<2�{]3^:l�)r˯�����>x��1:�b�홠M�����!�vwB^��]�l��*[����|;.�I��֯"g��d�d�t���C�6B���+6`��K�&6�c�$zL�k�r�U�)�O��vr[�Y�5�n�� ��hP�{�3S5��f��� ��ME�/%��Ԧ��ad� زh�V�S��w{���^}��.���o{T.,��fZ�z}	��4���0^VAh�=�x�P��'<xa$���Ĉ���(��7x�{��:��>����r�����E��;����7c�nI-{�wU�VJ�\I�̶Yg��� ��b����5z�c�!4��]4�0��=�"ā:R���?� Q���C�y֌,�`>mv�<��8��<O8��aOe۝�'���V� #�@A��YX�k�V��/�x��E�g�.5��c��N�-�m����i{?�e5��fs�u�Wv��R���gE�/L݈�˵��#s'�;/�ɜ=0���[m׉��׈I$�a�����P�\î�Nsq�)�'
 �n�Ͳ��՗)،p4"W.�������TH1/�o4��"r#*��P�Ǯ&���J�v�[9F��M�0�eWG���5�e��|S%�(D��+���$�86[��M�YH6�����; ڄ�w:Z��1i��#����?E�������ګ�w'ck�E�uܫfU]�����7��]`M�P�a�1Y)t��^��9v<1�Ou�X�I���U�N��Jp���ن�Ҝ>�[�G�u��|�+$<)m�մ�r[f!S�ڢ��gr�R�4ǣ��J��\�� 	��n�8B-	5Ԁptx��$�`�@�:�x���z��4=-R�"�8��<�	��"�Amm���#k-��?�T[���[�J"Q�H�kʴ4ϳ�W�PJ���á�B�5cV�ⱥ� ����N�=x�J\4F-��I�Xu.�SD�3c�p
t�x���:���U���ږ�n^5˱ܩ�Ɵ�A@j��*_8V���7�6�:c=y��a�T^_���e�:nNC�y��RcU��V����Zh^���vQ���k�ٹ�6�����5{��#(p��*sB47QMct�e�֨��U�X���BH�Ш�_��bv񍢿WI��lz8�
U;�U��<��)�sR��RÊ@��EΊ�gy�IqHP@q�%{d�0�f{V�-�a]0|}s��z�"�)��%XfD���ŭt�>���T�Xqn�rYs넦S
F�����aو�@z9�;��ك9Ӿ�:�' ۝������]���mY��z�a.��ᕂ���!?dp(a�$  9mg�ػ������S7�&���O�swū�����
�rk�7G^8)����egdjn�!�R��� e��6��{	*n���T��*[;a��ҡ�Yw��i�s�`��u�jd�Q�&�c�`��7�-��_oD�$0jZ�T��c��|�m�Y�����b�~�_tHJ���|n��+��LJ�r��Y���U�mk�mX���ki�O���P�t' ���Э�߫�o�@�}Kbȉ�QƬ5̎��d(¹&Qf:~���@R*h�&��0<���_��(�}8 �BK_T��h�`�7�ℎE���I�^�$����[�L�;z��K��0��m���%(i�|��p-���;�'�K<(b�Z�o�N7�X��#1��[|;��n��a�u�w����@{�(�N~X͞�P���@�4N��V1�J��9~���Қ��e������_0�X/�?6��@�$�cB��)�*ޜg?朷�3�\�=4u� ׀bA�����<�k�;�;��������{pc�_sY� �k_�r���66ê��,�<]�:X��ІéD����5Rĩ���
��sڭ;\�H�J&�K�L��W��MVia�-K�v�n���z۠c6�gK�߷��Z�$L)E�h�犭?e)؅� ��XJ��Z}
�id*!]�X��u��B��ی��u��(�6G��̈́��x/�q�b;#K_��w�Jn�O�i|���B�S�-.�9$�E��b��6W������[��H\���oܤ�&�?/K04c����/����g����p���'Z1�����l��X�z�]4g��i�"E�e��.\�F���5	H�F8z��X,�@!l�[R�=���s�	Ei(-�R�Q%w�DF	#{�����;N�o���.zW*�G�Ѷ����F4��|�L+I{~9�]:+���X!ɍ0.#9`�w��A�� �:b��~Q�Tb�'�&˵N�ab37��ՈA1r�����-�
��1|M�m��<	�'CY������r�0n�G$���'����� �3p0�䍘o8�"ym�t|�z��ڒwt�6�֌��m`�X
�B#R�����o�q�\�("��'@5�����W]�D��&��M��~�p���@��Y �<x� �b���c�65�6;ǭ�1�/T��Vm���	?�_���p���� �c�!�d�m�����
���$s)ys6Z�^��bOB�;�h�T��2�����M#�H�}�ո��}68`5M"<ȟHo�:}U��Dف�(�Qk�>��l��&���F�uë�:&��<��lh�W�a��1�/��c�Nm�߽��SW�[Mh�][�a'��ʩ��ȁn��)�K��@}���[�1���:o�2�/$ע�Y�Q\v��{��ԱӲ�?��IlJ��{1�̭��B�N<��=���{�����a37�k�6��fءֿ�����X4։S���N�C��FI����hT�	�u�o����k����S4�]'�Ǡ΄4��B(��%��򟭰,��%�7�`��t!��gC���[ U%����� *�sr�8�G�+W ��I��Ӡ���
`Лfz�Lg�_�U���*���P��cZnE`|#���D�J��1�+|�,Q��q9P�<��P叙����1��za��kTB�>�B��;���[rp�����B��zZ�|�K���y��a1�jhr��m�!ܕ�V ��?ϥ%�>�6���7]#xR�%���I~>+�X��驄 ~���/������1��^�K�?�g�2�xY �-<���N���G#�B�-�)��D�W��B�J$�39A3��a�vǭ�	��\��:��ė�9QFD��xcwHL)�^V��j=�?�Q�!Ɔ��/[;��L�J����|�,ٳ�ܼ 巑�}��S���$͛Y3nd!*$͡֐$�����|~rz��2lgMB�>f��9�� ���1��t�O�3������
ș
�5#���q�N��6[��P�πo���'�a�J3A��y- s���H{i�m,}��<�'Q��^	A[��G��LڈنrP�v�l�Wc����qx/6hd��=���1聱�v��[�{��4M(�1Ot�(�4pC�&=��ڐy���eʑKS�����([��U��Q��Qܖ66�K�㍄�龓�qA.�Qp-�+ơ>�xH���<��O���*�9��T���-�׬ #���1O2�TQ���F��q̤'m5|#|��
4��\��&�$�d�w������-:����l<�w��^��蓥�3���m9����_��I�^>=v��� >?gh���v�?�����G�Qబ��|��3s���7�jz�� L'��'�j�O�k���j��k�o�'fJ�)� ��*�̲֗�2t���/������}7�~��l��Y8�[��te�g6���Ͷ'��.��ܒ~�^.DGVkM�Ǫ���޴�־��}����Ж�L���$O�s3�)��Dɒ٩#��}�Q���݀�Qi~C!mc(�Zg�=)�霧Tq��p�c.!tDs'!<�m�c�I]�GI��R�j?�,~��h��<'����E(j��aƁPmu��7�����5��40R�vz\���S
]*����#��޶|��P4&��Q�'������Wݕy�2D�WjH�gɟpo����A�ΩL��j`��#����E�����П�^�֟{�U"����sR�g5���i�v�=��9��c`�ב$3������KĤ��,<O3&H�l�J�K`+u?Ŋ�m��>�b��ѢJr<ǗU�V�ʾd}���;���?�)uy�Y�L�G�Y�K4�k֓��K�EW�&�#d	�
ׯ�D�b��`�L�9���+�S����-_@}wk�b��)�� ���u���$�S����N�IcX��x�z�K��(� Ak����M q1'R{v�~'ș%>V bm�BY��jj����`�g��d�������k�[�̅5]0���Π���yw�P7u��oPX�$�S��ݱ)�f��5���I4�K� ��2�U�%a��[�!'q�2S��62�Ch	�"�_�!�Q�h�X��t��73�+�&Sп
��$���|�l��u�� {���:�A��G�8n�>-���m�۰�����@��eU��b���(�pz��c{ڰM�e�e�u�K��-�2c��}>��n3N6�,����n���)�o���=�� lwQ�хrZ��g�tY��#ג���a�å��SJ��h_�n�֚ފ�^nJ����Ac�Ͷ�)Lm��O�4c��Q-d*Dy\&
m��o@5SZ�diF׳g�x6����S��ݺ�(k	us��>�����J���	SKDBuwo��e���۷3��+R�b;�w�@D��a%)�pJ��$�u�_�x�j��pf��`uQ�Ϻ*g7;�~�fئD��ëFGW�F����۶�LQ�3����?�J��Z���<k�|���j!;S�ɜ'mȐ)�^���rgJ��J�oX*l�e���%�^U�daf��A�f��0v:���Hɜ�
�1�.MXC(���?Y�tmf��&&P�7����+�%�@�>m���;�4|��I����y� ��0W��R{k$�������<�+ Q��p3.3����M����]]��-_�G�hA�H�ɜER~[>�J�R�������R��HATۼf�N�Xj�=Ch���ޱbD��E�5�M�~�dDX�n��C�y�W�t��
(���>�q�ir
:6���-|������xt탬��0�s��D�|y�CWqV9�ߤY����p��z��[���AǷhFh �ʜ4
�q���u6i|��>�P�ǸU�_'��.f�S�� �f�����:{���	�����	_B��'�����N�ޤa�:��)̏��:�F`��Oe�2�=���܍4HZ0;A:hr��j+�OᎣ�����t! ���K�[������0`���ϛ����۵��]\�г��W�E�-�7r+���^��z�7�v[|�z>���5Q~XvA�xV}�b(4�x�j�#���5`�1�^6�0�  ��g�k��\�����.�Am�b��n9�0�ナ$	9|g=��n�s�6�����0�~*!�L�$ѵ�+y>(_ߧ���O.�BnҮ��Ʉ�$��]�na�9�F��3Zp�M�楤�X�zq��f��*�"ǼZ@V�;�&�8�:M��[('g�D.�ݾ��.��d���n�I,t�4ę������̫i3�ԅ��~�fզ[���8�]��>NH�f���ʾ��=Ky���� }�RZ��W�(qR�+DoB��*2�v���S���P�J�^���������'̂�{���	Ӆ��N���s����m8����1�J�W��ZĒ�`�R>�S8�0�sF���ɡ��V&_�)�#;��J�8=��}�G�����X��@ץx���������%�����

��y�|��J8%Z4\U-������g�P�+;�6�`@�5c�Զz5��}��$����ى`5S�K"f�Ԥfc{y/��F�H$�A'�AlV:��3����*�����ȏ�l�<^]it��	��T4�e�B���M�FDP�$-��:��q��K��-�[�#��,y�r�AbNW#�S��gL������X���_�[�q�k���|�5�	nG�l�oe��^�uihGR����F��.5E�?b<O�a��rUX�s������[?��9w��[��r3G����\뎟ػ[���*��g���C�j����R�?A�	7Y�O��"��S?'}6�] T[�OA�?��Q��os��Xk�*���q�d��r��]�۴{�+*������w�t�ogpeB��bwAE�w41.��4��T�H$u�y�5�k�&�v�e�~� �-`|G*~V:�t
�<����,RzZvF��DG�l��f{��ꅒ���N�$3FS6��hQ���snj�:Qǁš�I�ҳ��R	��v�.�_K��MF��6|��U#Y<��"r�7;�&�CbOIq�?A�M�i~�U�x�����ї��w��U��-�$���g�;��c\p���o](�.e^P��؟��Çe+󿊷GL;�~ՠ�&߹+��ϝ%Y5�jj�Jx618�sJs�
G�ȷk0����@�;�$���w�?r��&��� ��74u9�'��a�k�ZO��%���X�Z�|OnQ{ڋ�(�:��YMi:��Yٖ�WU�[��l�I��2FQ B�C;�T#��gXE�m���1T���a�|����T�ɕ�e =܃!��&`7�[����p)�T�/x�M��J��(�����LT��S��F�����p�ON�W{X�3�0�S��f��l)����EWi�Ei��\�'�N��"�V=NY/���	^N}����:�uAs���~p"��I[:T:j'���:��,��F{�X����F��Ɓ���D<h�[[׊�iq^�l����w�ח��b �F�A�f�N��߼k$C)�YKʮ4E[�~i:r�|ʭ����K��X�����
"��R�OT��P�j���PČB@���;u�N.�eO����E%o���e_2�B�}3tDd�y����>7?y��5ߺ䡘�^n�g���D��BF��z�����:�Uz�n�z<�׃, �B�H3�-*QZe���ms<-������f��KL<:/�T�{���;{jM��;<Uviا�(`^���n�=2 /g޳�C�a�����A8Ѽ�򏜘Q"M���S���}a���_��10�UP���*�=�aENn&�{U����`�I�Q���s5xI�@����c������*Ep�;��7�����4|)=����"'^�TΚ�̱^j��c��B��C�̄�����L�%�ф��H��{�9��`��>b�˛P�>K{L����y��^��lL<Bp�p��@g��Ńz���}��Di,��u
]��0T��d�����,�]�cP�_�"���|Ϣxh�8��I;�H�/pȍ�Ffo��>�2�����_��	��y��V<՟St�$p~��=��E���@����5Q�\^_�_��������_���������\y?�x��2�+���m���Pcl�.�����M��nr��D��;n)N|�S���W� � ����������!�m�OK���p�(�¶��������c8��7��U��_���C:�t;QO�"6Wz='C"2_�P7&�����tL�|��hH��V<��J�W��>e(t*m��A��������nzA>�n�%0t�r�����
��xҽxs�o��'���f?\�#�%*��g�G|s6�$�U��\�3���d���j���v������x��?�����-DK�o	I�<4�v��vX#����W�{�K$YuP�sZ5�{���+����}��\r��)p��~���R�s�Sg�ʋ�����r0X;Y PeY�7�]���o�K>�U���[�pl\��*�ᎀ~N{�|���R�.�Ɋ�*�{�4�F%�-�C�4�zz��5t���&	z�0l/��.e֘��O;����
LO��E.�ef�B/�Qj�9����B��[���8w�r+x���.�0O��s���CV����;�К���A3�H�/��[��r��+Cg��8FГ��r��l�k� ,64u�g�/���Hf�~��l ���JMWN�fX��p푋 DV��g�3��)KX�q�8���w���Ķ&Y��V�W�+:�I���[��%���*m����>ׇ��~N�+^�%"��pg�Z��u�����*e����M-�Ti������@�" ���#��Q�<�5��T_����X�}�I'���`Aq�N��+ca�97��������8�F5]U���c�����IH�сy�+��7����ATW��]�O��	ǜ�k�x�eX��䳜���xY)���LP(v��$ F�@���±z�P�����$T�7�������$縥��qf�vJ�k����<�}�ɛ��@�e'�gb��sG��@� v+�r;���l��{��������G��{�L����U�eApY�-}�_�n�Vh��2���Pm���4:bڊIR=
r�[�1��K�,�U֋l�i�n�%�j�,6�r�B"�+Q(+4QȮ�$Dcj�N�e.����.��B)�O����7�H����.=0¼ٍ�P�XU�>N,L�pQZj�0�	x�_`�5��ڲ��`� =Uc�P�����a�̃�{~�F�9z�m��O��G^�<t��{ɔ�`��U��D��KQ��u����=��Mpw���H�PS�����Ȓ\��:�߱V@R��Dm�5��s+�b�lΐRh�**irW���F����0h�9��JO#B+�*,����v�Y��ѕ.\p�X�~��a�#�� ��q�@�;����gV�e� ��rY��.-�Z����@T�ҨR
$�a)����:�x}���n�(a
fe��ړ<��%�*�VA���� �pb-h��k󾝲�e���տo��2v�c�.��״��{��r���0jY�m̵Jg�ܽ���mn�@�������L])�'9mx� �.��G#����DD�=�;����]�4gf��3dq�o��j��;q�==X�}�\�M!��t�O�&F�t�7���_z&�Ut>�=\���� �#K�ݑ߽���qg�L�R��ߡ�j�"sa)�	���P����g]�׊5���!H0�+�<)����x(���+
2��	��(�?��.�ZX>�����6	��s�"hmd�<Rp�s�4���雌%]l�oh':����L95������SLc�V�9�tzX�Z$W�V�?�:ѹM�9l�P�uE+���B|V1��<�O��.N7-��Z�cs;Ә2�w`�w*��#�	S�#�^H
�L��*%%]"��8m�g������]4�X�W"8���N�� �'�ާW�$��8�?�#����7Jey��Ԇ�V<,]�����g���b���q��ꈅ[9i0I�!#�����xOU`�e��X�Kt5�N
��6��R�X�̢�7���[�DjS�=����ۊX>.�y:��Y#�)�����;s�p�S�fz4��ď��Ҡ0��5ƭ�I�(-�.���,�<=�#�-�yn�-7���kĸu4��S�/�p,������26z��L�{)g0�Ǿ*�8���9�]ͭf|�gKwV����sxw�1�o�M���|�=�Sԙ��a�q��}��8Tm���{��d�]�Y#�S��t�à�w]K��HW���`�w��ԧnTc��]e�}�McV/j�-��+�P�S�4�F\��1ό�k�$*�Cr#���9�_Ŭ�J*�J�
.lF_��nB+�T'�2�M,{8|颭�e��En9mJ�]��M���3*�#=K�Jߒ>�}��|�(��`_�e5�$�?�^:.�x(b�:	���j,5e��y�
�Y��7�"y3��B7:���Oq��Nv����V���\�@DL����'8���
�X	��$<b������l!+���iyV1����sV[ S�^Bt�h|jV��5l�n �Ɋ�>�����׵��� ��K*��a���E"I�}���c��O�XmY��
Y4<�{Ƣ"��&]�tr�h@�nډ3�wQT���(.������1Rc��a�a�&u�� �����?G�/a��Kp�r~φ����`�(�v{BS��m*Oj����OJE�=��|��>W��9�I�;���n	��8U'6X�
��W��?��8rl�&\2qôd���m�,�8�> �z��CT�͚��gRp�{���s�lvf3H�V�/��lN���^9�FZz�on�(���fm�ɤ B�V�	tc�q&�{K�.Z�g��g��?ɤ�����d+��_� ���kX><��8�hֻ�@#^C��w�Z�Ԅ����)��>R4�8��������(g���wZO����=P��cc��ӂ`��Rr�O�,@���^�X(�{�i"�>1�9&G	��#첂�)��40�7��������&0*�ۨ�=���
2��H�g�[jt;4�Fa)_tV���9�t�ı;n������)���I�J���%.�O�'c� �ڒN2��&�p��g��ԨI��#Fn<x�\�����u#OlNB�{�n�KER��2U����tJ˟ʩ�'ʟ�!�&kÚbYW�z�楺����6��Xk�.2 wg������l�pm���D��@δ���#����g��JF�d��e|��g>�W�V(IJN|J_pG^�ߐB�gqx��3$���Ofy�M�I��?#~{�rn��>Q���b��a��9a;�hr��&FSȰ�,,[��g�]N�~+��K�Ϧ��Z�]��Q.�!��sO	Fti�y}��E��h��W��[0g�N�f�QU\ɊW���)ɐx%8�W�^EE/�qpeZ6�F���[8F��i�+��X��Q �|�_�dz��ڇ���rl�Q�{��;ٛ��˕k7p�}*i��٪P��[S�[����ؠu����<�B�'o^�'գ!j!��Y(-�`���Zz�Y�96�� �ۤ� �,���f�M�/�<)B���X�o�<�m�`�0���K\��T��{JE��wi>8<�:C�y�7���ͳ<�j�⃚mT��  ��<���t��Gb����O���ǯ���$+8�Ul��d�+��=����m�r��k��S�vҢ�6z��p�� ,���x3���Tl�1���-��k0\q|��Ґ�?򅭏��Ec�󏹑��������0�0�,���sZ�ue94I�]��ˣ�>��(�/�,���R�r;G�94��K��L�h8������A�Mlh��]�P#��CK�9���{����R��"�Æ���5Z�3Q0i�E��i�t�i��\�FmŎ:��w�[\��h����"讎	`?	�x���ZK�}����7Է��A9���Vg�DFwjωH�f����`����S�$�8R������g���:��C�#E�J[RY���.؃z۷qy�N-�9�����_	oO.߂��	sC$�`�k�Ӽ*i�6�����ﮞ���6�������\Sڈ�4S�����(�p1�Oԁ��k���8y��\w��z����&�,u����㷌}I�d0g1n��4�!���E^=��F��Z^�*qȑ���X�����:�������>7��n��TN��.����b������ҭ �<�E6²�P !�b&;�?�<��Θ5y�3�7� }����*EM~9�q�]0f�]U=�dQ��M�����	%�����<��n����%�m�c�{����_�懎���1�D�""l�	��;Tnqm��)�)���~� �.�r(ؾ�q
���GW{J�^��&�Q���� c���/����Ѱ� ��+�����m'B#�%k�ʙvwpS���z{���ʚ�̝����~�Kg�$���b����m��-8irȲ9;l�ٙ��3�Na� ]��cE[�9�0F���ݿ$D�'��I@��w��c�}�꧍�5@	�v��L�7����L@J�~��pKU\�V0#*����B��܀�C�9�CE�OhI�?Q�c��CyK��.|,Β�D�/(YWC�y����D����p1����"�#���V��
 w�&p�%3�!J��2���L�\-M[�y�=�Q���V���k5��A!�*z�0���a������ق"-Ջg��i���w���q�Ф�E:ҍ�/���E�1@�:+�^�*�"��oU�s2��k`��SD���I����Mu��C1�z�6��p���i�6����k��ԕ�^��[���M �#��Z��
��jՊ��y�r��t���BO}�C��[�TU�	�u+ ��dUƲK���J!����B���C�	��x]�v`x��n��'I��:N��xy��h���@<*ӻ�3�a�Ҥ[��������xM�Pc�C1�^�On��S������{�n�p��.d�\�{jZ:[�5�d�$�����:�8ӧ��s��K
m>x��J�]U�V��ANn�ʊ$�(K|��D���� �+CV������Q�.�lt�@�':~Ik�L�Y���G[s���R��{�藲�!��.O�~�=?��}Z:~�ś~=]��塱sJ�����+Th���^Ȧ��O�-��JO��ij�RDz�ή@�_�K�^a�d`�1I��M1����'W#m]NI0F��@s�+�0�% K�3���Ⱥь�M�m!����qI�5�n�q��e��Ͷ�����@<�F��v�t[�H��5�YVΞaI R��@���Vj�9;b���_�7uޑ\�GX~Q~�Y�J�G�O����V��깵����u
�T~"Q�a?'����
lॻd��Y�Q$�E)���G�4Ba�E:𥏎�d�G�SaE��pyj�G���w!�A/^�ؗ������]¶�/���+kh�cdrI�l�� �G�T�lA�n�ӜBAƶ]i���G+ ��*�&���B0LQ��,�>/��� ��FG_�֐������du|�0�s_�]퉓	\�)��Q}���D�����#۹��C���dSf�D�H9�� �t�������U�rXw�������eI�~�:UGi qR�e�Ni@'�cn�W��SL	�M,�#7?��,ZdÊE�f
�~+^�wf��������q0����5O_uf*���}1ֲ�h҇��/]q�
���M�dor\X�F����ՔbVA��!?d�B�/��$Z���+$����z|x��>�?�\���m׏�b�UpCr���]I��kB�����G�c%B��8b��Jg�^Cu��甈�@I�8�����,[�Wȷ~B��D��&\
�fW�xa����=�3�۫�y�(��/(�i��G��d[0�S-͊Sم�ĭKȈ���0�Ц�f��c0n�]��-u�:��R �3��\oeD�N��!Y�~/yݐɭ��P�n����K�'��S�D ��,TQkJ��g^�Bsq{,:��1�;',�n��k2i8�/�I�|��M��8JM`��>���Ͷ@��q���$J����#���.i�Mn<���ILaP�_���6T�zA�Cxeb[�������+e�`H�Y��8���V\(��q�����K[0�9��A���uҭ���� ����U�ްGxu6u(�@�T��R���?�be�����5	m"v-0ַ�p�e�7�C7�ʉ� qZ����P&�����ŀ�v�s�67���!����4 l�]�yI�թ-��1G�P'|�|,��p�C�s$��%R��OU��A��@$mK*z^��+@�:��k�G�7)�Z}�3V���������5��5�5����(W���*�c�>�I��L��� �EC<�e�7�r#��>�����L�ĵ�d���I;���m2����Q7e� y	!k�܊x�Y	���T��e@��G��.��$�|5�Ws����f�G�j2�u�H��}֮��0N#�D8,�qO�\' ��(���jM�<$'�i[�ub6J7��@G��ig<#�8�ީ��EjlI	�~(�q�_W�m#h��,ck��1_³k�����V�yc�����<X�JF_*%٩��]��c����½�U�z�����j��l^�sf���EA�D�S<?�憘���ˡ;r`Je�/���%ޯ�M�t9mz���� u&?�r=�8��C��="�����a�y��,�3�T�ؾ �I4���j����)�d��K��,p�cOR��콶�� c�[��_�7n�D=�=E����
��7P�o�A4T����l��veit�js5��D��,RZp	i�ܰsیⰁ��.p���5��>�mfq'��y���;�j�M��+�5�-0��$� b�۞���$�������^��o��i�2!$�Aj,�J�ۗ��%Me�p(2�� "�Kc�.I y,��b�����w����8�+��X��2�2ێ +�1?WǸ���q+`q�l�on�o��@5bJ�q�Y�|J����o(_ì.��Y;�?L��1 ?� :�!��f�A�:��VU3v�S>���/����f�1b�I*<���n�Qg`QWqP�-��yAv�Dد0�������@�k���JN��ЧhBZ@0�H��cd�)!�]4&�e��~��W�[D �O=��	�u�0������W���[s��}�f��$�h��.h�qV��>d��\vlߏ��w��(8-���b�D�o��F޼��b�	� '6��V�,���o<�8'7li~��u�ߡ	����2Q��4��=^:�ga��xU^.�]*���?��Dt&ǉ@�
RJ�?7l��.��jpYX��gS���f�z|��̈́���3���X�Y���'j]�@���>��ծ����F0?�[2�{6܄��\{����G�p1�I���h�\hy�Ka��m!����gV�/��v:��k{{m�q.Z��h�z�zvK�&��������J��ņvŎ
�N�<|6���4ݺ�{V�.�Pf����2D�֩l3��cŧ�5��0>aħ������]	���O5e�;�E*U�(��\��9�,F���;ń�I^�掮�~��3S���L���ˆ&�<kaF[�����1�{��l�@��p�~������m���*�n�m�M�Jv{�	l��}J����L)����@X�]�~u�u1�u}�)@��]R�Q~.�;�p(�iC�n皎걟����8�G[���25���T��y�]��uy�V|W�`M��)-�]L����.U���%�Q�U��/!ĿSߝ*>o�z�~/��{������q��x����/1(b�s�PV�h�T�gBY)�E���k�����I�DG��U!���z���a��}kf�"�h�.a�Όe��(����/�L�����=�y�+�����ӳ_�� 3X�C���?(`�&OB|<#�h�q��g~���'?�����<��%�L�OzE� ��6��I�����D��G����4�~}�\&ȇ��!��ʶ�}�E	���RlԀR҇���dбI�~�
񏻞3�{�Z۔J�/�Ϧ�V�t���w��^����X�l���I��'�$y֒��L��DT��s˱�g�L;��h����E��,e;�7iU\�������.ܳщT@�l|R�8ڱ.�ywS(*8^�|X+Dv{ɴ{P�͟� ��:�#���F�6�˂�9��7�;��0��C_[�z���*;!x�$�/HZ�|/?"{����0�#��~'�_Ekb~�]Rx���
�E��c�S�#�*�5^`z B%�'|�"���̡�����v�F�Ŵtc����Sl����6���ƅ>OB�PUcK��x��zmz9h�bb	QҡT�	�"���4��t'yO�ZV�g����#��oU��2�i�5��l�
B�+rȵ7h��:�HV��R����E(�r�,����e��Gy���q���{TV�ngb�����7 �|��4�C���h��=�;��M�n�x��i�N��rvs��Ƴ;B���1�*H�\��?�qb��FY��T���t$� jl���Mj��
�Q����j C�/��ý/�k��uQY�� �2�# �b8-=F�7F�pE����\+<Lj¾�M�WC�N2Rq����Ϛ��Ųn���m�h��a>c��E�)�����D�2����*�� 
�ޥ���l��*0hSV(��Ed&��YG(z��G�UR���L��`��3����G%" ���:�.���<zb�P�q5�p��EX��v��~��F��D�DEh��ݨ,ʩ��ľ(��UJ]�Bhh��<�Dy�:��r�V�؎�_�,@꠺|e^b��jĽ��NԄ��/����iU9j@�pl�����5(�������\��2�\Ц~��$*S[�&:G���\��&�7|�%�֒<�޻����}gsD��BxpO6	�6��oT;���\݀wC���� ��u�xD��gI,�Rg���T�� $ĉz�4��e���>�#U�H3���G/��R�I�_�~Q�Ҹ�p�w�޻V;�h�J�	�c��cu�E�&Z�bAz9G0����z-�utf18E��fc�@%iU)7�7Y�n��05�n�|Y��%V��]�&9o���:�>E�����b{��a]�6H���2�ym�4���Ӈ�f����sgꁉ_����d�vJM��Ǥ�'}�����jJ�g�\���[K�u��b�V`������Iy%�ژ1E�v�/��D zT��hY������h�xB��W��졍ν����?@�����a�A}�6�*����<K|���1Gr�P�Cg��#�7�^��]?s	A�aG�������DT�mi;������K� _���0��'
|��7�C<���uӗ=�v���Ζ��JDWh>��KT���j�uNQ��N�Xႇ�/aNCv�:& �k��>ƹһ.� �ϩ���p��D硩���.Q���`^��u$�����U�8�{�BC��t��x��6R<���]m7��,��+�BwI�0��1���Ԅ�~|���Z�?�ѧ�Z�wE/wߊ�f%c�8��]��G�K2�_��k=�.�K���'_�H��B:U�Z$�$:�#��R]݊���iU�$��oӰ�߾20�6�`:?�Ue�TTi��r�����d���bH\�Ʈ=<
jq����K@�R���V�dL%Nd��
�'�n���p/B��'M-'��a��{3aɘ������o���Et,0��������?AO�XC-T���6�WT�S�����Ao�Ԁ�A��/m<�ʯ��ĲfP+��4?��ꜵ�OV�B�!��Z#-yK�>��uP	�4��w#�3:��?	���sk-��v�g8�V�Z�ٍY�m�m��[��r�\*�?a4����[& �	(�v�u,�!}O$�I>���\JL~�ha�n���eh`^��Tn�C}��ՒqV�iezO�����z�����ݔӟ%�;z���,�Z�DG��+����C��%.?8��j���B���jNl��ǻ��9j�"�1�@��P���ف�����;�kS ���[P9�o���T)_���+���X��%Q�xT@`{/xA?��+p�����g��F���2�2$���5�	m`*��Ec S���#�s�W�*7~t���ȼJK4�dp���;9_�X����@���Ӗd�-�����Y��nn�p�/51X!�wN3�+A�ΰ��������1��QCo�ijl�9�LCZ�`�-�
��\<�˩z~==c�4E�)3:�2�E�?s���ؠl�֯^W<v۞��n�2u�^c��$�N��^2[��ٗG�K)0�xݐ����e���UI�#-7�=���
���Α��@"$}�{?�`��ᴖ��P%�8��ڌ�kD'���|ο:���[{g�C���U��~)\f�W1�$��-�*u�~�����b�E;z�e��2��,����z;���O�d�G8�Fl҃w�������|`�� Ҡ�[2~����۸�y<�*!�z�2��c�Ksf]�m�s�$�S��b:y&��8����Rp�9�'R?�"V����U�����g���񘉉��`��V�\m�7�LW���f�5@�\,N[���[�$Mߤ�'�9�athF����?҉���-�x�b��D���K.�%P�dK�L7�����'x�`f��Ԋ'���9I�Wdb���a������^���8R�K% �Hp��y~���=S�����̳��6ߙ�=T�7ڷUKtF��p����	�����~W&f��m�p]\Iw�5 �>&DMU�yleh11����������G��'{V�Iɺ�S����?Y�ʹ�f��l���#<���G��x���a{�R��������e�L�72��)��#^X�6z]��,��rq�;f�D/�C(��ҙ�)MHHTƼL�8�dV�n��zv�&c����ouJ�.cS��h�o��y���]_�C���f@�8��~�{����!�������F�H� 3�=!k� �"�S��{=9�9�����2�:-K��'�33XD�&_KÉ��f��л��Z9P�� =B44~�{�����	-'�k1�Y׹q� ���I���xc3����$�#�D1��H�{� �PbwO�x>�o�G's`�H�o�r�n��0;r���t�����Ȑ�s̑��nIu4�oѮ	/*o�Cqu�W�B�עJ����\�y@�Q؀Tgg�>�2��Ɨz��<�Zv�ó�P$2�~���'qL$;S��4Y�� +wk�p�h�����YE_����C#Tw���Ha��h�$!��1���VB�8�z���ڝ=X����bc+�'uG��N4�6S��O�ˏ���J���[<kN��o��@�c��PTg������o�*��09!i
�:5�HL˟�w/�٣�ߌ��(
���ȡ�\3O_MYP�D��,�E�*�v��D��.g��U�hUH�%S)�\~Q�D�N!���J��g�}A��Oh��2Y�=��4y�����~�(}(sխE��XM��Z� �o;m��	?��ޘƞ1�x2Q�Z�OLl�8� ռap�U�=�}�:8�d9t���dD��� �H�Ȟ��SőȰ�J����e/{f��H��r�E�������[��N�,X���}��t������J�N���Z�;��Lam�t���1o�q��������^��r���jO��2��%K��Z��#��pR����D ]����Cg��u��-��e��Jl��K���S�HFU�i��Mr�0�!:Ȧ�{���O3̞�i�𮌧�X<�8t��q���a}����8�<�n%��=������A,%�����Xe}Y��K�}�^<U�����e�a��f��8J����(XX�	k�v�o�|��͖)��6���)�8�lᨂw�Mզ̀0�F�[&+}O3u$�c�v%f�j�h���5�^��E�,�ZY���d��X_�&�N܎�)1&vF��T�$W�F��%�A�iϝ��g��$80 ��o���c�iR�ߗ��sq/w�\ @��a�U�M�dKǐ��d��e�ހt�6�{M�QH!�T����k�O�?�I`��)�r�+Z��8]߅i���lЭ���[E;�
�.�� ��<	�z��f`��T\�^��#�}ɝlf9E��#�����?5�C�M�cð�݆�ϧ~�j@�ϵZ���j�`?Wt�W'-*ɷO*_0��'�#gΧ�c���OY;�鳇�)� �]�fY�N�F�Җ�޷��s�a��P�"������ˈ_C�B�n"8A��J�񧐃�B��0���� ,�e�U�}Yn�:�\��Z�:s�(����PR:'yZ������7gbI�W������@ ��F "�(�j���k�[CݮSo��'�1��G�Gt������a/
` g�36�`򋵅Q��D�*��
j�8��Z��x��Պ��C�bW����cVc���@W������O�L�!r���Q�xkv�����QZ~PԵ�:�BG��M֓�wE��=�y��3$7v�\��Vq���H,	�0$�[U�NU�\{2~	���5�_��g^.��ߒ�ɊU�s_70���4�C$�p>[Ð�K�#�"!叆��g�X�9	�.a<�v8:�}M�H�����0����U9`�Ow��r�9�8qwFg�b3�`�F�R�`_�^kx�@��p���Q��K���Z�Ԋ:X��~����/`c#g�ylr%^#����V�!L���}���e|��O�ׂ�V!W����-g�t�z3�#ibEr�+����Q�N����d��^���KV����s�I��`��A�"������ӄ�ax��8a��D��
��~���:HX8|�Ɍ8O+�t�{P����5�$��/��a�R�����O���΀Ľȫc��Ǉ�yL?�㍣Y,�{�=[�&��X(�t�{�#����#����P�5�k��9���Wh��鵨%hx��9�K8��k�kXDU��op�@����:T�������9B#�ht�ۓ&�~��[s�<�C�jYqKJ���D��� ���$uV*�8�@��0���I�g��-+�S�/��{k֔�;�����Z~���N�{��\�%ó0ҟq�˷��~**D��C���o�����j�H��*��4:��!��|��M���yFS"���R�ȉ�̷�8��c|����R���VoL0�z��g��S�S2(;���H쫰s�/{^]O�?k�������72�z��_�cx���pLD���rK��Z�c���W�\��<�~�-'���FE� �;FD^Cx�gڑ|3��m�����^��X)�?a�[=��B�5��A�]��-1�*�;u_b?���H�N=��`�J#[��U����B@��M1`�[]Nl��U�IJ�E�� Hlp6fR(�����mnk"t��*X�����K�BzDJJ��h'���$8��@��5�r�������Y�L�=��	�uҚm�u�����!C����m����iCoV�Y���A���O�����'��}^��D�JLx�����-W
�04��_%�\}_O���IG��tYX'�^�n6ᅏA��B���G�rH���K��v~w1�a��\���:VOe�>�f%n���	��9*��CR:Y[\~�]�o�b��8	^�>	A������f���#	�_�\�_�{��}�ȕbb����R�acƢ�Xŉ�T�Bqnɚ��_]���vkU��s�Vb��h��D�p�N�\)ǲ��`� p�21}�+������56����H���#�Z���ʈ�ꤸ07GXg-�(���0����,�������I��
ѐ9������~UI���~�p���������g	L����q�:�?G�$A�k�+�%v�M�d�&�=5�R�
O�E�\A�C.��_��d���RNn�����mu��1)V]�~����o��GqF�h������py��/$�0��ǩ�Lv�κH�׋7;j��{��|F�xoFl�r�d��^�|�a*!�{�?9�0������Z	�'ڲ����:/F��G��u����wX�de�d���T�@ޙ��k�6���E��"�K����h�yP5bn��|���&����Y��T�2�{�R������w��:UYfN�nPEa®VT����t:�~��ʫ�~����4-��̷r3�k;�g�AG����Viý���Ӂ�e�6-G���XsЀ��ڬ�UV�-O��J��ϱ��l�����W�E�Q��.=��X���i��3<�[���~A�
��y��w�y�_5Y���?@s��$k�#�Պ��c�7(̬A�-}��|g�-j*V�&F���{`��j~\O��#0j�+H�#VȫmԴ�ZbP���[#����2��{������B�o����^�9�D��rEP4�L9���]��gꎥ�e���)���&>T��(�:?"�D�ǭ�(�����^OwR�zߊY����X��m�M7�:,[i���)�ʗO��\EZ��S�42A=�� ��F@G5����C�se	�Ǧ��}bc1�z_,%lAhM	^b$�®�ң��~d��K1{ho���qO?� �ФytYx���W�w�u}{��9e"�c��������(f3�7 ����B18AM���������	(zם��(ـ��jv�/+'.}�ab���!1x{F *$�<V$��Vky��7����+|�M�9/��J �ܴ΂�����
M������~p����Z����$'�J��	N�t����\%�%�Z 2�f������le���RP���ϊ�Sa��*0%nfu�)n7�Kd�Ԛ-�v@�Kg�;L�HV�E>D��g��E�#:1|�p5E?h��&6�N4���ؐD�.�V�6D$Oއg����\K$�� Ͱ��n��8��p��w��hz���a�m�ȍg��HB���Z�a�����c��hy�&�nJ�{j1z1���4x3�9Ÿ��8W����	'Xf��Z$�쬑�S)��<�����<rrF&I�����֞3 �5HU�O�uC%�Rs��f-"fUP-JyI\���O�'�]\[�@l�6����@���iM'V*�;�,�K��":m-`D�6da���P4��wq��L�H ��E�K!�����SR�~Z�ۨ�ڿ2��u�VA�]z���?�����J7��u�F�s$c�t)�MК�����8���%�� ����'�r6`*%$w3o������[h"� A�G7� ��	r�%�^<��~����'��Zc�F�p��<�:|hӌw�4"�;�f�w6�c�4."������	!�Z��TUݚި��׀nO�]x�{�u���5�p��>����i��U���a;�[��I��oQ��$��%M���&��|�"� �]����p�C �G~��m�C�ϒ.�0U����\��wb��fň��ߤ,[,^i�}���D`k�%:��̤��a=���Ig<��(�j�Zx�9�wIm&A�<�����p^l��ށ/� ��^a������R �j�f����n�o�d�N���%��+Ө�7 ����d��Ƃ8!��ĄF�jD��<ZM�ʆp�F�O���õ?����_���>XA��ٙ�q�D1h�L5uJ������N;�	�u�
�9=/� ,i�P7a�o4�V0�$w��;׮��2�u���xDF*㣦Ă0Nd�]1�}DHm�p@��lV�6%���M�n��䤵=Px$�ń#�d��8Ԟ�S�p;D��Az!~3ZB=� Ώ$j;�G�i��&mn�mt��i~(@H��'� ���W��hD�㲐ڜ��k�i1���o[=����Ҧ' �|O2����2�d��(E�]��@�f�q(���lhP��9��V|�׏��5a-?�XP{b:�#$|����zUO�0� �Tw�D�F�$Z��'���9L�ܳ� �Cu\�����<_S��THW���}�1��7�`b4�4��g�Q�,H%�`���Ή���)�r����eU}�vL�X?�������+}*��ΜE�L���Z%�5#�	C�O�N���3�v�^�$�"�Q�k�d��;iX8��S�����E)c/�"��/��H�n�{��~�7k)�x�si�_j#���2ܨ���������s�{���&�)���Il����Q���cһ��-z?!�����	z��F|��å$	f ��:��y�R���/,��	E��u�(�V�l�S�����h0p�2(�;9by%��j)��w��C�)�j���ٴ�T�3)�^��V�P�f��W  *9�\���s�p�.x�3]���:!K1c2<v��V,R� ��
�A�+�6�0n�O�E��ɫ�����'F�=�M������;p���L��A� �]'�f�����.YԨ���~���%��c���V�X�Lo@���H�����z"#��W��xj�ɬ�/�oP��k[��}D4A��Q�cLoE���9�*HA�(���:���I��]�����/�%7�.�rr�*&<^ks������%��XʡSg�}��LB���04e%��I-q���2��Q����Т�ڱ���r�w̲ni5��%(��j,Φ�bz��LV�QXvj(�$U|���+aWF�̩fYtr+���a$���m��|F`V��"��nCr�>�+�_�������1�}�%څ�8nՂ���	Dp���Wz���[��1��MTۂk�?�\�.
� �Iǵ ��%9�zފ�*�^���D���Z�	��6;��޶��买+�3݃��D���W���G�J�
��pp��?|Ǚ�6�/?1��O�������F4���� E����Akz�m�X���[z�?R5����h�୨��N��(Eʝ�lYm-Y�}A��UC�JF��W�pC��c0.���e�9��t{+��5q�OJ! Ys�'���X@�5�x�12֘��>����+�[8����NC�����tcv$O��LK���*��\\�k�;mD�Dӎb���=�I:��{E��k��2�NZ�nf~\z����/��M�i�9v��u;ґJ�;���s�(J*u'r|1�=�d�K�cG�Մ�&�7����@~E�eF#��cĄi�`��O3��d���B'Y����%��^ZbHG�f3�c,�^��e<�HBT�}�<�n% ��y����,���sQ\f^��:V�g/MC97~��;X𖉻/��ڣ<2d���=��
/�*,i��̈rcb�NI��OT�Λ)�ʌ��*���δLò�C��?Q�r�����b�&N"�Ш���P���@���v7F��-�g/�V��^�e�wlI����}w��w�xǇ��Z� Z��H�W�����u� E��~�[`a�D���-�ˠ�6F���n;I���=�s�z�Tn��u��ɥ�^n���Y�Sؽ�a���bx�H���Y�����}�'y�@m�|����5���2̒n�ٙ��n��'r�^7	=��������g׸���,���4�̉���I�ϑ�Dپ165Y�w=��%�"LG{�M2�:5�O��iE�K	��Д�Yʖ��/�j*c�±�*q¤vw%�h[��/�E8d�m` �E~������6П�ͽb��sn�RƍZa���,&�3KiLGE�I5��	.�7\Q�:S*����}��w]-}y�C�K]	�	�ٽ��n�*8�P	�0��4"9��\'�����	VJ~�|C��������/�B�O
>��❝@L��U�ޱ��Xp{N�	U��5����<iQ��9}XF���C���j��"�4tm|ص��e��Lw��F����HU�Ͷ)�L�y���5]a�o��)B��'�!���.�˹���HNk��גE1r���ĵ��N�F^�'c<24 ����T�O�a��cw��L�h%Ҙ���W����[I)"��J������.x7��J���i�/'YXȈ,�Z+� yXm�ۻ�@���z�@�-)�>��"���D�i��Df�m(�F���?�|�L��
�7�v�Zخ��349�8OR/0���]/��\KP��\�gу�K�^�כ�'{�%�ʚ=  1EN`^����(��Z���tk�z�4����c0��A<��_ǟ��2��`$�}*d)��'�Ӫ�	�Q�Zi\|7h�(m��:l���iz��p$	��K��r���'7D�
hOg���r��v͢� =v҄�s��k��e겄�8���)�c�yS7�!��Ƥ9��)p�� �=$(��Żۗ��y<��}	��ܵZ}��۲�x�Z�� �)�_ĬД�S'D�q�Ķ�L�&�Ä��5��>?f�� {�PM$"��*�T�:��` �U���!!BZᅘ����E�iѭ�f�Mr4>fg$;JS����sz]�+�w>�0 ��	{S�f ��Z9�9hq��j�q��пْ$sX5ұ?{�O�(�$���&,�ѲJ�C�ކ�=H��R0�`�5h���%TX#Li�������S<;�b�n����Cm%<(~b2��5�'�Vu�䙼�(��̂���"�,�����ցz��W��"RmV�3&Z����siE[۔�Cހ�/�(�G}���[2	������$�T٫��X
ev�BR&S`�����b��$���@���9��:��ʜ�����X�7r�[�l�x16'��E�LL�x�>�IIy�_���w�awF�2��"S�p�R�펮��Oλ��,��`ӎ;r!U(��tԄ��En晹��9��*�ޮ����HXɁ�]�����C��@�:8�\���@>mK��ؖ>;B[@׬��s�����k|�BE�Y=N܁�d�!tb���DW��Z��i|?�E�[5I�����%���k�S9s`�u�u2"�x��NKX����/�ǀa���#h�������Ąg��D���z��fO��<@������b�D�Ҿ�c�x/�B�:����%G]��!P|2�T\�/ �
��$����o�e�N�J
��&}��Z!��CcJ���Z.��]Kc�d��5����c3t�mts�Ȣ�_Ͷ��9.V?�%��˦���J�3,�u�V_���W�rX%�d��.��&)#bߪu!=B����I�qW�&a�����̳�ņ�.�m^��Ny���p�HW���蹃�����ݗ�2v���\N�z���.����	�}3U4�=�GFq�M����u[�S�C� �� ��J`P�A&��`]�]B�Q�)G�VIw>���I�**x�I]��}q1����m��wh�nbGm'�D�."3�#�L������Y�M,��|���)�A��-��iա�����s�Y���Ժ��-��#��Z����r��!�X�|U����1=�ѐL����ӷ��q�LaŤ�3�=�+l ���d6_��R�)�,�#�F̨nN
�F��[�U��ހF�6dy��߲�~����;%J���{$�g�(ǘ�E��#l�]i��4� {���J���kX���l�!�mt�n��;m��}�=
|v?O�Qմ��I�
�l.|�<�4w,&
n�p�"�\�T"k��4��鹓ڔ?�>���^T��G����k1o�^�%㰣��(Д�ٽ�E9=�:����A/t�2�|�Ea���ܥ7�7r����%�̚p�?֍��}3�Ca����c�X[u�{n�kQ��l��������u�S(_V�9�K C�U��� '�9�,���0��G��倡��Ξ~	Hɟ}��{,J�%B�+էЦg�/Pb����0�#]�r�âh)�}֖�U �Q{z���d�䛡ਏ�% H�{B�
���V�3�H�Ð��:��h&�-J� Em�\:��
o6�9�0�g%ȫ��"1�8����M15~�������.�#ZO- /����d t?u�úZ�Յ!�$�b�L��4ۑYX�]���;ia͂	�r*���Q�S�'H��M�j`��uNq���:��(QH�5湀�4�9*Ґ坫�Y�YnQ�&ѕ�s;�r���krylQ����Y�a4nBĥF(�Te]�n�2�b��~�u{
Ӟ�6�n��Y'�͜xd# �)t�1��ۉ*����K����j*�*�����c���F�ilL}�Y"�]g��\%Y����xA	X+�"����d&q1� �I�.��|[p	Zn�w��?�Za��w�_3�#V�`[��swH�tُX�r7Ŕ{H$��M�{H/zW.����P���M��5���q��U�U�
`�$��3��v�>5T>���V���W���3��y�E�9�L���y��d�c�	�|�2�)��6%?�XG�R�Կ�ލ��ŉ[ťd�0*�!]����Ӻ_�>��n�Eӫ�L���.����,���:=`�|S�H#$��� Cz�6!�RF�¡�׸5�>�I������2��,S���e�4�j�b6�W�^?Waq�b�w�tf�/8�[�k%\�#z|��aW�Lj\G�i/Y
��<��/t��4,���4.�R"�.��(���T�o�A֤}�kuE�h)t�mVĊ��(�ו�K���3���+��xk)�@Q�H���w�0���6�d�BY�Ǌ��w�nA���L��x Y�H��ٴxҽ��Zֈ�������]�s#��j3��K���$�=����'(@\�� ��4��3�:I��5Nr��= T��a�&�ō9s{�R����K<����+�8����	z�<��x�yވ4�EK�K��EVNP�D �wh���*<*Q��M��;��s�����j��oď���#6D�v	J鮸F�RF����$t�~�o�v�V%*��U��/��֮Ҁ�_�O�2��S�� 2�h��m��0t Z�5��s�om.���L���&�)c�<�UF;�x�y.�p7���n��r�#�n�p�P0-J�/�m��F0��0Y���X2�8[�_K��QN�8	�AD�-y��@��=Y�e��(Z��\��h�Έ ;�F=����~4�/G<K2M���n�u4��&��l�?�*"W�W�'��I��V&�	~�n��v �J�]�?�<ܻ�`���C��un�d*��p7�ewҵĎ�Nk&_V$ب��D��,��.�� ���O�qN�"֣���X��Wp`�6���>�bS��*���>��4˜c����j�?�W�/��=�9#��D�v�_���!�a�+,e�D���R�C����D��sR���x�F��rE�!��� )5�!�RA]o`J?(�;�ih͚B�����:v����h�s��&ל}�h�i�Yq�t+�{�cΏ��k���h���Y�!�5��q���o�T���=��t�5%�?]7�V0��DfR�s�I�n�K{Ʋ�v�S�Ku�p��Z�rP@w��� �˶ʉ1קQ�$c!�:�	�X�QS��q���1	�t?F�ޟg%:0��;X�:��ݞB�rw���e`���R0��gE'�0��������Ǡ��;�$� 秧���lo�7����A��t9��؜��d2��l��gh��������r?�+{��X�2?��ͱ{^y���K���×���+��̺�����R'�q�Dv�u�+�z��,�R�̴}ޚL���RZ�M�(�[L����>O��m��+ڵnR�u��e�JYB��۳�L,�#�))��!\��F��������iK�.�s�H�`�Lo��Ǎ��⑹���]b����	Tވ�jl?̄?����ҕ�Pv<�G���g��A�r��Ҵ�k��Ω�]{�֓�	 �CO��"�x�8�J&o��~?_��j[��/�}̭��x����?���W��O�������j�*�������5��y����ID+Y�%[ ie2� ����h°Ȥ�sk�=8~��Y�_�N<iCp���*�/����%�P{����U5O����3�t����W9���cs�DM	׀����}��c��H�k��p{f)���-BڐC���Iyd��3
�ˁ�<y���Ѫ%�J��
�'W��=�L�׈��}s�oH� ��,HA/��[�R|Ha�����t6?3�ź��g��1�+3}ѧЀƙ��.s��^�����8v�Ւ�<0�}U3T$O}ڡH�7�����}/�Ň* C)����&w�|[�	��25�d�P~�����%G�7s�����*��*�������.��`�L
BE�㛉�p����l�-Z�_�����Iݶ�4�=j��n޻W��h	=��Do���s��v���)�.7n<��>��H�?��
Yl�#��ۤ��V��B�K���5|K���^��?C�(�+�XK��U���w��:�\���myȻ<�4_q�4�m4��@2�rߝ��|�Q���o���T���1K(hz�	�`�XY����ޡD�$&�Ǐ�L����EJ�e�X�`�Tl��n��cL���v!�x���n7� (�d��y_k3S m����!~�*�[Kg  X�b���ϗ%�ˊ��=�>�ck,���;�
J�PG�C/'0��^�>�MS�?{mբ�a�����I� gh�3%kEi>w�������}���M/kLɑ&$���U��K��&]NG�mA@�����:���NR�k���b��a��E�:G
B�V�������s2VP,1P��O�*�:g�g�!��:�na�/�U�YkD�쬷0�|x}�tO���I�Țw�B�7������zɞQf��s���^ ��!�G!-l��m�$ic+��m���Ky�(sÕ��@�z`c"�O.9����Bt�//L�3]9�R��ǔx�w��?�+Z���a��3lS��29[L�QݭZ=�B�	�Gf?**L�wDYvy��2�Bh�#�H���#�9��N�5�F}2q��t�����=7����;$1�E_Br��@$��m�� /@ �Y� ]P&�	r<	K�=��B/@�ß�kτ�3�p+Ti�C��K��"Zm�c߄�M8��[tO�m&�+�~ԂFm�� G9��R�t:�C%td8(4���Տ\���l�NS|H��+�!�ɷ�U? �B{�+�QB:)���P�p��pw1�#m]���D_��&`�v8Sf�(;IbI�8���v�.κ��7DI�����L���sU�Ig�m��j{�)�� ��1g�ԩ�����Ԋ�||}W�c�ʵ��%o�H������v��<K.���~�<�LK��s�q`��f�Sd��*�Wʙ�ʱ<ÏWL\�I3/N`mm��N�p0(o6�'E�u�+�B����R�9*9/�!��5���ؗ0�f���ǟ�x��^ ���� �'>��~��9��uH��W��˥����5:��8JժZk�L�eQ���ǯ����F;�(Τz�/����[`�IC�p�8Oa1,Y��R��n/�ec�1�(�aUR2)@��F���P�K��@oW8؋�}웅�U�k]\fS�;{\�6#@jv�C����ŧ��
zsA�wX���/�ƷD@�s��Kܮ?�w-��ik�4��0�6��"�\���+:{��[�-�E��4�~�N���kb|�@��f�D[�ϵ�(�l�0�8d��
7�۪��po��vM����m���c�S��������M#��dƼ<�V;2.T�|���7X`Ԣ�  ӄ2(�Rч��R�o�a{�3�|�@� i�N�����Ï/�r�����/,�旆*gG/�is�p��
r��o�@�z�)�l��<>XgV����_���������; K�7�bۻ1Z;��7��O_#*��*U���`~�nn�� AI�K����^�a31αS)$f�H�썗_��Z0`��Z��o.'�]�O��bX(N�.����a�q��P��B��.���j��+��Nb���Q�,)7m�Bp����X -�(ٶGbG=�B���r?�cmV�����n�2���\�0�X$�קe��y�����#S�`��$�B�3�&8�(��P�j(pG�G�����!b�Ʋ�M) c�����L������C\C�ʞA�3PG��%O�^Q��B�S��BqY�@�/lOI����5�p�'I��z,��#�I��p���Z�+�p,]��}l�c��k�,D������ί\�!�6[�#�h+e�o4��C�L0{�#�|D�]x���ȼWT�`�� u��^yJ�/���x
�~;�3"^�=cg������5Ş�ٴOw�t�\/�x�YAR�gȱ����v_Ϊ��*>�m��~�i������خ�n�g.�qq�-��҅f�3����#�M�����!%�B��sT�z'�E�	���_�[N٣��G>���Y7Z.��KU�Rn������<ǃ�$������aQ��=��1/�	�=�����x�Q��o��1?���<�K5/�4���]d�l�̞k:��?�$��@���bķzui��}#5^�p��$4���W'
����WM1`0X�-��L5�[b�Ǫ{/@*�T��������ty���cB9��?������R����Hʁ��&<�>��'�v}���ɿ-1����{Ebf�>$�Ǟ���*?�H�@�V	��8�}�쿿��TQ�Q��]-	)R�Qq���CW�9�7e��xM������8'����� �*���!��z=y�� �W�*Og�H��TR¨_�h��﹘Q1V�1�����W��]���^%��W^�Eɐs�5�$s{��|2�,z�ua�¦yh�iUM4Ź2���f<9�
C���u�gh�Ia{�B��}qI<�y���'��d��}D%��{�f0f3�܄j.\e�uW�!�Z�M\/����'�\��^���,G��&�[P!�2������N���v��h�\fq��\?Q�|�m4�5�\������M"\���̪J����b�kf�����������s�r 8�	EP�`�`�����F��da���M��C�9���k�)P�?�g48H8���X��`*Lƭ�e)z6e������cjM���_�-$�::4.�)(��u,=κ�4��[�%�MkK*�mG�»�.�~�8*"�V��-6�es?��ʦ�PNEdu�vFH�]_]�k�CWT��{�h����h�G�I@���������gD�����bB��זnx#�'�� X�]�L�[<	0S�6�S��.�<�T���n������� ����.4Kdt�n�sɘH���N�J��@\C@���r��E����0�S��Q�:�$�l�
ٶ�r5��60�'��Thr��k�U�bz�@���>��k7ss]M5�q��fbc�"K?^��/�S�=��?A�u?��j�V�e��qj�/������)�k�����q�o���J���fZ"������V����/YR���=}�P�wei�9���w��;���6I V�u��eoq#g���i1N�=��bw� �᪮�""?j���)�Եr?@Y:Ůn}?
O���(�AS��ݴ�x�nK�il� �+�7GbIz�]K"p����� �o�8c�M��,cS`]#ͅST�z�IM��Jb;@���+=�.�{���_P"�~��L��V�[�[mx�JgiC����-K����,���+$v����.��i��[�l��"`����H��^-���o�n�I=H��eIg�Wnfz�'�҅<YA��Aj��âJ�3�UVh���]�����Į��M<�_P����Y��!��w`o8�P���2���C�j��}N�����EYxsR���n`�yΰL�	�k��v���/-�5��u����T�����z7��+8�L!Ĺ#�˵kcL�?}��c�֩[h��[O��Ø������^O�m>Ө?ed(:�h��}�Оt�(�DU��.��k��ϟw	m��^��zܫ�f'i�2f�4�2J�[��d2nW,��)�lݝ�����KNq^<�{��kU����N�����@m�����$���Zi���wHX�bɆ�ꗷæ˦����]���:�2�+���QECH�۳N[�)���z�-��if�D�M00����[�?K�-~�4�	�9�7 ۺ����Vp&�_D�m��� x�[�}�N�n���ʼQZ�9�7�1��H��m���b5"*�z(�a���e�N��+󉄪��I�V����B���ɶ�!Nwhɪ�iao��Q�.[_Id�vdL!�(@G����3���W,}��x��q{�x����ϳ�jā��qآh%s`.���*�d�Yqym�ɔ ��������4zQ;"���S>Hg̶O�M����{Y���p����J��2���!1�Bn&Ʌ\�gΡVB���"����Pb��cB;{�Z�T��<l�pQc_��3h�a_l&�gw�s��w�7W�!<��;h�uz-����F��[Of!��E�7%��<z.�1�n��i�V�������3��	��D���JI
�u��PVI�/ĕV�
�>`��;گ?,aZ���TUN:�/��K��[�F �5�j�)��|�6u�{4�����4c+��D*�gD�E;���ݪ���A]�/;fe�m�h(qz:?܊�*f/�������|p�G���^Ql��\�G22Aʎϸ�>~G� k�nsyӜ�Nd��仄t��zMުٕ�K�>2�lcN�[�:�>��G/�}g�O$8f��H{��Ѽzv^������*>x�6�a\J&��n�Q�sd��޵����/��n��I�#�>c��o1�<�<��piz�p�hJ���R�!�-<���X)����xg,�ʞ��D#�Eɯ	d��.�Mi-\Nh���q��=@�S�xL«�g�X����]wj��k(P��Cߙ�����^�Y����7�i��L� ��e���q��-S�����r�0��J�#���c^�w��i�"ʑ1����`
�yj�s� �k��[����x
�M�.�ʊ�vP�`��Ci�����_�����9Os�3ƾ����FOkg�:��T�&��X�F��Eˬ,�I<����O`��~?��&p!3.7�L��V�����D�{]�������6�W�?����7`Y^�����HABEt���
��1		�u��{ +JN�n�W���0tAjB�b�������C����ŲR^w�x�ظ�,dR;�A��{5P�,@f�-nՍ�)ώ�B�e�^�}�C�l�dG*��C׾����M��׳�6xμ����O��]I�*�s��a�����I�nt����.��`�s2?���{�l n�d��A��i��0g�vM�s�\i�$
R.EVm�Kp#l[Tt�k�3���Х4���m�il�$��"�/�ã�����_�02-ۈ��M������~EE�t���۟p�/"�ۜHb����<�_:6`i"��^�I!�/����)�4K���2"����n�`=(��mگ��e9��	K�7�)�:����^ ݦݲ aW��#��*��1�/S*�[\��}���2E	���I�����s��i7���@��-#��TE�)K�G����U�b���{�!yUq�9���{�<	�yo1˥��Q��q���[��]�|i������_�������ѱ{�������^ X����5��g����C��Q4��\�O�"�ͮ������ӂ���)H �*U�i���EfH�u�<�m�� )if��*m̤��c�p������&�f�ܡ�Bə�+�O����_[>�V�+���gF]�R8��� +MA.�/�k�x��*��O%�~�H!��	H�+�Uܠ�w���t5������b�I%�Ijv�*��Tf�)	P)PZ�}��o!8p����b�ﷆo�/1p�V�nN�1T�b� �PB���q �t����V�pɽj���t >��~�ƈ�l�]����%%+nj"I�J�od�Y���cl�	��7&er����=SKʰ�/�yL��d/�-��(�� }	������N��U�s��ω�s���B���Jظ|>���� =�8�1o��p�j�S�}���L�;�(�{z +����v��Aٞ��s�󯓛�n&t�od���j'O��v��Ύ~I$|�_2�j�ޔ�
�4�2<8~�5ؗ�c�$���8	�و������%Q�k��.V/-����ң����-F5\6���T�I�����8C���d�C��sA��	���XV�B�n����u���jt�0-0� �1�dR	,���tN���'�k���I	z%Ϋ'V6��L٨#라<rk�r�~�3u���C�q���k���?�A��־L`��Q���9��ϝ^�W����u
�O��u��rJ$4��8E\ܫ�қ�ZoveB{���BĊE;*D7"��-��º�w�mb_XERnI�Z�wS1��M����vW�FF�Y���L�6���t�����¬y<.������I��m�[�t��>o�4����_���q�q�*�C/��J�7ߋ��Vf$�ݾ����~\�I�W̤�
�F���o�6���h ��Rhf�	2�3,���J�+���1�e

\���|j��J_d:�������<g�[��,>�f(wІ��O�dPXr�ke�]�[�,�ӥ
q���r�E�ž7-��o����oK�t��EF��'p}X)'v��8�R��b����ǰZ�٩KC�aH�6�q��5_�O�3���iP1�z�TVG�ǻĔ�}�j�|)�w��X�D���t�4�H��1G0%&5��Ä �ƭ>��2�x�̬��*���'��ZVa���8>�ħ1�&`X_��8��`K�aꪮ�D8��7֫�[��W�*���l��yU�O��q����,�R˨޹f6Z�2�E�c����E�M*C�Ó6NT��IP�B���?�m�i�������w��2dNJ_&��O�UՕ��ެN]����p|Ӟ^ �z�p�蟃 ,S��L��s�xoaHń�{�,Hak������|U��e@�s���gI���tX Q6�n�4�6G�u�l�yՉ;
z�'
Ǉ�wuޭzPw�_� ��p���Y \�U2�!���`������� ���(����v&�?�
��;�hv>�fI��F����9�dkrs^��o�$��!e�9E��,�	��O�l���L[�wp*Q�(�"!�3�=�B��>�E��'�#��_'�kچ~G)�ug����{���dl' �w,�G��Q�x�
E��|r܍�u��q��(��U���;i�>mi�e� �5㳙|�9�0��8��Ġ/~���;�����\T��$-nY�q�4��p� �;So�G$��T�io�7ꊲҧ��0�K�\�R���g=���&�a�t:cˬ�Д�����R��@�����Yt��T�Zh�fO�C@�ʘ�	���p0�>yh)Dw D`�5}}1�ࡴ��j��n�wc�aY��RE�ct�>k��µ�>�J!�D�*}���]cTx7��m{���4a��|:���O�8HZw��[)1�����o�⏳e,��O�#xG���"Ե�2=��x��� 4
zɃ�C"���b���tP��B��/L�h�^��h� kv��S���#�8t�'!❇q���rh�@�as�pfm?�?�zM�iF/����8�l��ӓ���T�ݿ�4�}�Q����|U��N��栨s���O����ȑk�4�%�T+T�O����b����X?��r�0�D���5�̷�^�h�	'&�1j��^�h�QC��հ��JQ��K�M����M׈
���&��3�{l��"Q��0ٶX����=Y�(я0u�J�MUY�G����j���嫤�8�E1�?*��"͘�m�!��l��E��|E|[o����x`t�/�79/�m5�9;�?.%���������������ƞ�*���p��_-w-J��G�p��Q�lO�`�p�<lM��_ub$��L�t_��#�3��'Q��Z<e�q�����?K�j����`��[J�5L������Z��VFk�g0^�n%o��iìx�LkE�������:���:N7����+������]���hs9c�pND �j�9�'���a�*@�B'��2���SL���}�#�Ţ���\="�p�q���m�F�z�alS��&�H�E���J������z����bp�5+Q��c��Ν\9>*gqU�S�Yd��n��Q������:vu�����?���"�\�'�\�>���\�L�
*�!3g�=x&�ZΓ:�
-�'F����x�@���ӷN�%���1����޲��I���
�6���@�M'�F�?)�k����%��?�kJ�Ջ���&�fH�t��ұ�z��g8�f,�e��k�	�S���/��UG���l�-�kwע2qe���ۦ�Q� H<� ��g��#F������?wc�i�\�0�&W���M���-Zfʄ�b2B���>�x�2�/�jOX;j\w@m�u����D	l�p|��sm8�'�r��q���7?:0g�)�S�l9�߭�} U���W\{h�P"i{�P�P���b�!��poFD�3��K�&H�'�>>?N��
�|�z�����ʭ;Ǳ���>�Tɂ��&ܲ�c�D�IM���ل~�RwJbWa��{�GBo�H,VWu0�1�<�spJd��y���U&��İ g6穲�i��qXp8�$�{��/{�x$����(��S�ܘ���:Z�C�! ���W��°s	�JAb���܍ɬsuec��uTӫ�c$���՝Rjl�F��@�е��`���6�coj�᥮�璍��$�ð|\����܍�& 30����j?@$6;�,�Y�Ŵ����9�������x��` P����՗��Jؚ:DV�����	:~o���U�_Ҵ�~%w;���BG���>p�y�M�T��A�!:�T%�WKU�p����!�4���%��-��C���5iZcG���Y��/�| 	'g!���V4#2�6���~��#`����or�='F����ݞw!�Q�G�ڬ��%S4.�]��5���{��.�5�&k� ]�8��G6q�^��}d7"P���P~a}5y��x�)%�֡!%D�%�(���P�a����@�E�q� �`�)��D���&���x�A ���)�M˃�Ô���۲�� -W~湄%=7�8��"0,/'��y�V��ǗS\,��b�ۆ��Ě��`f\���e��,[�?r+<)ӣ�pߙ��nBi�Aբ� 	&W&>6���@��(N���zQ��}����=��sZ����Ψ?�F^�;~���}�R���mL�	#h��M��1�-�v���n�F/��k��	���E��٬ٝ۷��(�@������3.B�����c�5��z)�﹃.ĐB�!/�#4e4��oêb*ıa�*;}PF����`���b�'et�3�ـ�E�T	�9�?��h�H�jߔSEy�9	s�1��U��2i�Ӊ]L�,M���y�Z:�WK�r �)P=��ԝT��K�Lm�6��mi����S�$�ϋV�Z(��[��]Qy%K8�k���������8��M�Tt��x6��b
v����.+�d8}�|��ba�z�r_W�hu�;Ӆ�늷9D&�M�S�p+��˝�st�_8D�>A�R���Q��{雈 ,��������2�h�����F[�9�w�ͨ2���~S�~f�)Hp���	<(1N�P��U� �?m��6w>��JW(7
w�¯d)�k,�7�(Z0��J�"dV���0��]vَn�2��F�:��I�P�R�`�<G���ܟ�������
�[ߠjN�����<���<�f��_M��g�ӗ�`��LU�ǐ ��1�X*ze��ׅ��H6�s���~��72.z�<J#��(Ѝyz�X(�q�
7��	������n�[��ob͋pG�̓��[ڞ�Yz�0�VA@ L�&
�/�C�S��"�d����/O��:(.�\��������3 �?�q��|h��;}?�7
`���QAŔ��[dT�˜K��<�Ƥ��Xɿ�i+�9d��Q�me^`
���Ӿ)�"��F��^�#�u&4����G���M�� Ɉ��~���m�vC(���}�ԫ�� �o��<Eg�� �CB�*��WS���3�����19a��B�$�#]t��@J�����c�?E�Q��jӝڅ4��ܙIc�!���f�x �H��'<q�d�5c�*bYh���"G�M%����e���b���h�~C���	��I�Mr�J��uab}�5���z������iT+�Dm�|$���_�Gi!%z2Q�N���ے��S�	+�+�JJp��B.`���-UGM���"�%(���n�i;����V[���(�K��ꆕ��A$4�Օ4Zg;)B��Mf��iM�D�R��h_x����6�J�rjw
�ui!�{Ơ��\������R%]��h���c��b�g�#���=5�Z��N\}Xe��*M��e5�G�cnpz���t��Q&T���pgA����������[�
}iejJ�P_|R�x[XZ2��xI3�9�E��Z�i������\������q�v�¡��xT�Q������juyL�k��
�6���q�g�����N���4���-��]��c��Mz�%f�/W#��Eπ����>0�EV;��6�#���7_�?�B�T�4H%�W�Z�cY8`{b���kC��s���~2c]�}��R�f��L����t �b�,�뵾,G�x��F>&�JYx�����KW#���N_��i�p �'��=�kFsz7C�Y�Tؕ��.���Nc+m���iz,����7��-m���5-�~D�׬--�b�/��� ��ësضye�
�g_=�:����A!��jD�ꎮx�,�j,��u���T4�O��Y{��K�n��"��P�n�_J�u�P���5���15�!I��ڦ|�U�De=�"��Ȳ5�\H�J���������o����{JD0��E!��R��A���~���D�%xnNؑf'ETdm̎�	 �S�~�O�?��{&jK����3� ��bHB�1K��:4IT�i�~�w� z��~MƠ��n��|+/��L�����u�_�ͣI���P�UwYE_�R��u���_(e|���-.�w�i����X��)&�jU$qU����:Q'�n���'�%�򌭊���o��PƘ_�F� hXQ��Ȑ���B���Bh����26{]u5�^+��c�^0򸸴���q���Jy�P��!����B;S��;����2��mDѴ]z�@o�lX�æ�g��o|���b9:擌�v�h�{;�xzpq�gS�I��ғ6�s�Rz~�D�_;��/ñ�m�A{����<��4�9�>@����ފ��G% �c�=��E�otZ�K�C�.w���<C�Ρ`!\��w�HG�b��[^��݀�= D��gdiԵ�V����dPcqDp�/P1���0s��3v�5VRA6`H�ޫ�T.��Z_I3���[O�������dyJ��D4�8_��Y��c�T��<m����ar��;&E�FT����ܭ�=3��H I)�R�9�;�����K���z޵������/�\�^������,{؈����g_�}�f@�g;�eJ�ຯ��{�������V�M���g��`q�EY�)�>^p���벭�F��c۾<�c�g4!w7<����ceªǓ�7��0��	�&H��J���nF�p3�9O�0^`E�tIs��y=�.���0��}g}~d+�N;?�q�2 ��@x��Bd��H�P��d�.s��o����������r�&�"��~`̣�[7e��C ��3����^7p}��~kV�+]O��;z//?b���5g̉-Ps]�׺����~��c")趲��lH"�y�U�:���]�Z��J~Hu��G9{z���gu�ӹ��[����QB@�@�8�"i�����U@"��2��6ʤ&h�S�r�1���)�.�~� �_8�^�є:��Hu�A�1��g�r���v� �	����fzy-����ǵ�1��%��+k�>������~�!�(h�4�1�p°�&�B�^�=�Dز/:WU0��3x�c��D�`��a����A��1IR%��P�? C����u
�\��=��Z���l���X�������5/������m�6���DD!M�tF�ut[��͠��}�vl�Q�!�jtr	�`d�Cu�Z]�=�s	!�J�{'?�J>Φ�s
�;�����l�;�����h�1�cT�o�������6�Ч�g9�P��JӦ�0}50�k�P/�D��Y�-�n� �˰Y�c�Ǯ�ʑ�)-|S{�>�x�0��Dt*=�{pM ��} {�����BKW��\m���r���O��&�eI*�����3!ox{�73�Â\mi��Rβ "䀻vs�Y����vEi�A���U�+H����E�|<�v���� �U�Y-	�XU���&�ؚ�b獵�oU���*�S�iH�r,~�#�v		yK�Җ��*e�����L�U��-E*�x�#)��+Q�2J�@��!d"�,kb�gq*��̚'^��4��a�Ǌnɤʂ�`�Z54\B.d����#M�&�L9�I�X��1���Ȭ0Y��o��W�ШڄT���;�>$.4��W���G��.�	�&.N_�Z2q?�TZ�j�
jC~+���Z雂EO�E�#��jR[�\�)���c�����Ԥ\�n�ځ��d+�^�
�ψHfD�Wvt�]�0e��bȒ <5����LS	������A��72�r��zە[��6�n���?��Á)��.���=ķB&-*�m�1�`ѫK�j�K��&Z��y��,��[�� E�C*�>-��;kϘ�ޙ�.�R�#����,L��c{j�kt��'����X����d>׷@7�E�S�h��k`�DS�Y�]����d���cn��B�">S�T8l��|�q8[Sj��w�s���)K��.�M��ZM�[A
��J�K��/��ֆ\-X`�[�D���a�:��N��/b�=dE:(�����s�C(>fϺ��bOX��ų��볥+�z0Z�
��x�x]F������6s�Jdlu��9��9|�6K���3����� -�ȄrblY�8mQ	��I9�Iu"���f�Yl)���ݥh�b�����yWଧŲ����)�Q�EZ4������an9Tv����(�-�6��7��ι��D��D�T�bq������%���_�#�x޶-{b�n�GJ����6M_v���}��`(�w�,�o���7�α�����g�c|�����|����/j���:�1#��#j�>�:��P.��#o�7�GX�/6��Oa�.G�C��c����ݱ��"n��TZ}Fv�5f��10�t��+<Kn��%v���}Z��X�I�,���Cc���<w�H����Z��S����!�wiu ����XD�(��&���g���J��.%�B�j)��Xt���x��X�~:	��s��ʐ5����;y���ھ�
���.O%��s��?چ���Ify7�X�a�ˍ��!���v�,#p �ʱ0��/��񁉚<P)�OYu`�0o��h�8E(��Mʇ�4�>���tTˌm�"�F�7��K�<�j����� �v���C=�����xL>C���m^`+D���|Zɏ��+�x��-ot��Ay<	9����]��r�	��qA���O0 ���	��������Uc��I�,T��o�L|N�l�.����XP��`@M����u:ɳ�O@!5Ku�?IƵ�f�(�*�ѠI���U���l�L���;Y_�P�1)��O#������	l��<�d:h��ꔻdLD*�A$P��o�5C�Rp|`4����ġ�P�d��5
C>q~�,����*���^�S�M�llD�-O�T1���Ꮌ4�����N��F��v��*�p�P�d+�r�OWJ��O@�F���5�0h[b�}�Ց
�L�c�Wz�[s�t��G��>U7����6�x6��ޮ���!S�r���{u Ѽ��~����+��������}K�}��i0��L���Yd�%���#T�GhmX��������?ռ����	/�`n���r�vQ�<�^�Nܚs����k�4pdj:�_� d��|�l��u��#'8�T�C��տB'elX��
Q��|FdJ������6A�[Ծ߇?:���9��\��RX>���$<|^:���7����"x��󺪄̏�	�Z6=s�77�X�/��=j���������n�Ϝַ{�D�E��.�ۈ ]�.���|�X;�L�C-Ǹ��ǋ�C�a� �&y��p�*ߢ}�Ո�W*-�r4Q`�k
�;}�/���)؎������'ocv<m����i��#G9!L_(֣�t�-gȻ�P�@z�ɇj8��b���P͘A ^m���������ۍ����i�	}�uo��`���T�>�\�`'�4�h�oCJ~U�O��iх����n�/�J/y�]�)��Dz�^/a�\�Ɛ��O�=�w(�f���ov�Đ�ߓ�,�P�\��WQE����<�CU�u�V��f�Z��1u��8��θy��T�"��@TkSpk��|�����T�Ho�Bb�a{���f3-�o/��{������V�+�M[5n.<����~QBѮ��.Z��@��&����=��>��c^���/���|z��9n�D��0DgH�j78Z�5Y� ׽6aL �����W� �K��3��&8�A�e8%�"Ff���4yF5L���"�Zk�=Y��5Ў��Og6��:C�},�^:�i�c�E�|����seKڱi<��׎�G�z�%���1�g��o�k��a$��jD���d�1�_���/��(��اOېf�y�'x�$��k�Pd�$�`�N3kJ���d��%�T���wp/��UZ�'؝*˓%Q k�m�� �����W�s7��	�5��i_6�R�pkbpǂ%ߢ�1fь[e�z �g+MM�9��N��*��Fm��\��q��+$��ɩ�Ƈ`0i1�~U��7B�s#��]a���1�F����7Uh|���ÿyǿ
6!�����%���U�|�H����MS�>}yT�A�����sL)�� j�u)�?d3��C�/RW~EM\�t���~�m9�>x�`�:�N�c���I�ZV������S˅N��ϐ��Y���`���b�������T,���f!�g\(9\v��&��nC:mX������]ZW�et*�'263��\k�ag������Jt~������)��u{Bm7����hS,�`���H_�:0\�����>��A��ŏ�L���Zя��g�x��d_�:�e�d�͢��N4�J�z��	�?@C~yt0Y[<5�:��:s����	�Ġrq�1f^L�q5�+`�������N����# ���r1�.~3*8���(8ׇ��8y�Pw�z�o�c�5�:�����(Ʉ§���(��v�����%8咆���8��@�5��_�X�5����>t=^08/4��D�\���k7F&� nG�M�h8���A9ǒrJI\IL��)�ru՟�ÀIN���p��*3Q���0l�=/*V�s*s��A��Ǧ��v����N�Jh�I����s�ZoFL�P����Um�n��BJ�s�J����I9���$7�;)��?<���NaP�!�(%W`�t�4$z!2������>9.H�
�a3��2�S��]W%5�Z�v��ĳ�kp�X������Վ���޸ �o�f�p,J����'�L��Zat�p\�UZY/�ˋ�J  ��nU��3�](,Zp&r�7�jʓ��l��V^�{�I-�F�v�#���R�u�پ���w�Ǻ������/�+OQ���5 -�IN~Ԁ�R����e;�	i�"��a.�CAzKY=`!��p娜�9�v�tAk����M����W�;�k��OY�nʣ�
���S���_!AC�G��	��T��ld�w5��5v���9�pnİ1�/��u#����VPh���P��˓�!��(�Us�7ME,S�����&i)i'7@���sv0��u)�t����Yu���K;|���6g�	VR�0HG�M��	.���m��n�QNmi����:��=�P&�)ؠ���T�ڒ�V���?\���X����IvP�tg����9��8g]�ӸJ&#^1k�Nd��
8Z��c��
��P�sI�� �̂��嵯��IݳYI�㗟��9m��05�\y;s�=|���_�	�����%�J�T�
�~B�姸�cxK���JE6��k�G�=��Ta��'�jx�_.�ܱ�f�����X�b_�:t:o��V���M�ajĽ$�&�D1yg#�~���^���uxe$�x	-��-�����([ʃ�e�KQ�hj�ʭ�c��Q&�+�����Qԧg�H=�`` ���4@"��i[2������V+�8�܁]�gI�� �z)��3䈺�"[�E�^U 3�>��m0%���?�\¾?)����@���Ŧ[�?��c�6�!c2B��ND�V;W:G[��O�{r����^�7l�^s*�O23��:�g��x¿ٝY�|#9���W"�cn8 S������˝���@�迕t�&��xIJF�~�{q}����]&%V�-M�!b��J_��)�V}������9�,�TR���� ^D���)	��{���ڂ��H=\�C I�[[5%1aPU��U�W����L@����S�B$��J�q�{����fT)�G��&g��;�l��:{f��sl0�1e��M�U'F��۫`'L�	������
HTF\M��ɿ����o�U�D�s8�z?�2�ܙ�y[��Z/�7�R1�iM���S���E<��"m'��|�:�A���)0������+�R�����G�"��5�q���*Wd��p�׿���|��!��۬[����� /K�$����λezw鸾���P���ZA�D|$�6G|�W1���U����&^J��{��������� X���Kr�� ���o���!�Fˇ�2ZnZ�W4��N�6��A�{�v�J�z����+�mly�gM�,߈�uӉP	5+'��O����<�`�6l�8�A\q��=,S�I���'��dꥣ{� K�y#Ty��FH�no�ϣ(�[6nK/r5�^vC8@wg���~��eb��p4a��tK�lO[���U��E��؟JǱ�A#y�Qָ�rZ	�U�k��`�c<��T��9����B�[B'h��S܏�w#8Yؔ�ߓ�Z��ǲ<}.���1�|�i�ӟlא.�8=
�ktֶ�����}�~�����P��3��|��`1�mi"����-2lÈ?:��h�U4�t�ْt� C�B���������. /6��K��*�a�Q�ަ��)eA�^�����C�Լ@��Xa(���������s�����{�f=x��P$�G����
��&H.I�l2��YU��1I��� SQ��݂NX��y\�P5��oɊ��k���c.�M��FՑ��~be�V�j='Hb0F/Y�F��Z+i�a�\==�vؼ��Ao��~�[�I��|�KBg���4�C�=��������|E����r;�RYp��+M;t���Dߦu~���[J@{\#�򳇴;��]��p�C�!�! X����+���h�4#�YQԷ�%�6�̋�[����Vm�I��_3fM�n�0T��r}}�CBd��#Ү�\�aT������?�b�����xn=���Q����IT�h�����	�������V��ot	������r1Y3�(����y �B�)w]o���� 9�GeBNցH�N����X>f������]��kB�)F��cV3Vȷ�NHi)A{Tm����H�l�0�,�ƥŷ�7�8w���k�]lw�O9��H�[h$_�~��޲��aC��B�q���g�{Ǆ�oB�~�#��^�p��G+%���^�H�x�|6r�E����}���O���'?���;	$��g[�k�I��ޥB&�O<�a�/fhpN�Bq�>Hhv?�D���i��mS������[�Q�4<��,~��S�V�5[��X#j�bv"n�l�� �܈##쩗����>�Vm���=�x�Yv(h� (�)�3@_�����kK�퓱�ͪ��Q�I��߄�=�hQ�\�9o��V�kq4(`*�o�_��&��g@�NkE���~�̍�;V�x���[�
��G°s��~T��c��\(�:"�2)h�R(6ʸ_SϘq�ٽ��{�g�1.C`J���*"�:Ҋ×�ax�2����H�b�z�NV?	P◤d�F��c�|�'�&`a��G/y�'%��zs�' �+��?��~�;��-ƞ�S/�jhnpA��fZ�,ˣiG����	綖�͡�e+4߸w��C>�������ͻ0ޥ0Y���RZ�H8>���5P��V�Aj_a��n�f��	�$S��t ��D{W�������5ڱ�z�S64A���12H�n���0�&����8\:]�����%���5� ��db���V�!|�N.�{a���kr�hpۨ�U�A���ĳ�2��WB k��c�`�N���}����t���M�l̞��oԴ��B�e��Qv���3��0c���������Q�m�%1)��=W�LX��T����ʿ��K�rt1"ʗ���1*?��^#�A��F��u�t&1�{�1���
��� ��O30y�H�ai��|��o7� ��%��S�F���mL�S�|B_!g
����W,4�noX:x:9��_s�Z/<W����|4��0�I�>/�M�jB�z�~��+"��K��������1G����dk9��>�f�̼�#��G�H�,�?R�e��f�@�ʋ�� �N�a�L
^m���%�v7	F�>��#$y����;�D�~)Z�|Nݗ�6Er���K���.@m����n�Хr�[k��6��?��f���Z4�4g�c�JU͌��q;�ɸ2�����fk3���߂�3��f�w�)�jZ?�o�r�P�'T�h�?�2L'�S7/b[؆�3L#��B/6{�����OH��+Q{�p{䋁n��$*02��j$j�b��q��e���Gp������H��\�#7"�oC�#@k��
q j�Y��Bz�P��V}'����ّЉ����6�Gu�UeRFfP��n+q�Q�_@��5�4	�Tg>� ��M����2�'d�I�L� ,��dHvߜ�����-3S��$��b1 �D3�wo��뙁#b"�H0{�G�*6f- �ӻ�O�4�z�;�sF�Z��_j6�п�"O�%��,&���#>�T<g�����mx�{6/�!ӫ�K%�Lh�ѵ/��\~^�h�\U�]�R�Н1��B�ᜏla����˗A��롪��o*�8��=���V��K:�,ȴ����$��rDZ$p �**���[1������j�@��h�*"�-l~�֌<Z�K��b�/$��h�^��b�R^X|��	W������ ��3h�!z(����3|���U�gF�	�ǗY-j�rL�s�!1�diza��?!����/���$���F�%�Í-iIm�/6��Rm�ň:�Yͨ����C%
P�Uވ�b��\��fÁ�Qq10�D�KuWҠ&��vոC�{�����M�H��f��|�;Y�:71����12���4#U�R�^W��J���+y��9� L��19�qw��������8D�\A\X�{���T�뎄��m��*��v���a�� L��9B�G
��2�T6w#���#��]&
�nb���)\�CN^�%8��2>jO�ZH��P��g��7����A����g)mOAo�j��AW]KPX�MC�;���M�ۏ��M�α}�~�w��%��nO��E�$��[)�ȳ[�~�=3r���9���RK��
�G�;��$�?8�%�7���)g���<���<�a�䄜��$ː����N��j�H/b�Yl��r��a���B��+W�j�)���:��$�6�aޠͩU�(�	�6t5솗k�y"<U6cثnO1\3>[�<Q�JV��]��@ߙ|�N{7��[�Mm$� 
���0Ȣ?s��������-��-%�+�8�t���M<5�N��m�RLe38oa�?$(4:B�znA.�H�6����٦.6��Y�ᇖ��ݡ�J��=#^�J��V`�Ax��G���5����	���K.����5jt�3?ռ�E�2D��!�)&_�%�vΉ�rBuu?6���Č͔�\J �ٰ�)^4�w����oIe�΃�i3μ���0f��$ɤQ`��3(Tv���Xx�+�����5�,3��߸M��d�1���� ��b�}IU^^X��<��~Y5[ݦ�8�U�r��i�p&�)S�`X&�dB�����mk;�s���*Aڠ�A9ד
����8y{R��ʲ���m�7��qy�e�
k��F�Vcv�4��1��[5D�Co,�c|Ϙ<WGe��0�X��/]�'�i��1�͕�����N(��
������_���i���Z�	j��"g�Xxd��Qߩ�p�Db�:�1�_�GE��9�� ɹ,���?`t5�飵�aƦ#�C;6~zZ�Oć�-�m-��;�C��a�W9���.ۓNX��nU��'�%8�8��j�LTO��.�a�!h@_�5p��>J�i���	#%$�d�a�ItN�dH�	j�2D)�[n#c��*�}`$R/��&��:�蒘[���#[�E�l����UY�fr�娝�;깭���*��nɌ���P_|�u�3g3e�O�%׮�T{l�zzg@ӽ8VY���̗�S姄�@ʹ�Ob/\�LES�fI��
�Wȇ.壺+��}�5ƣ�]O1�F$���r�C6(��3�v7���M���=�^!�)�j��Ȑ�#D,���8����Y a���DзH}�"����~�y��cX�H�/_���n��kq�I�(r%PG��� �uOq�������)����J�/-�����v���2��r�0�5��0��g�r����>���OtG�f�̰[�z7����V]���dw��bjw�Յ�WK���[q���=�	�g j��E�U}g"��ȡ�d}�c�"@3$��xU��V�]m$pਜ���E�q$H�e�NȻ�$��{`�s~����h�������w�nQ���B�'ЦY5�����}�p!�4{k|׈@p��<���]BQ��͉c(�L��Er$�ְ��B$����Wf��ͺ�K�����[/�)-R��aRb�4��G�3�S���n8K�u���$���!���q���,��]ʡoŪ/{^z]<�%��wǰI�b�g ���/��ӱ����o	�o���� 6�ْ[��5�`o3�Ǻ�����
h�,Z�����ʹ�U�ֱr_L�O�W�!�h^"�k!���O��'C!�/�D��k�o�,,��eZ#/v��[����N�1���]pK�E���s����hƇK�},��iiD�?4EOu�O��w� (>f�8��^d*��+ACg��x[ XRE�[-�}�]0�jM�SX���v����O���)N砄
 D1N���צ�k�os�I�Î��s��4�I��d-��4�Q�J�
wCݿV}��E*�bЍ��Ța�fՅ\p�R�7���/v��)rE�K#D�%)���Ùƹg���d���y.TK��٣��Y�_����6��:f�*�㣫	��A1i��+8���?�M�׽��E�9�4��)�.A���.6`,���ZNR��)�M�ۊf�"[GK+�9}��<g�y`s�-Dq53�?�tt!��yҔ��*u�T�a�_�+��关�5>p<E����_�aQ�����aXj:�8W��SC�G,x[ȊS��N��;��Xf&@��8�Ũ�$��D����3{�wGI����%2�=v^78r~��LA�Vy_h��߹Z�����_Sہ�Ԫ�p|l�WY���XJ����NQ!�����^P����ݢ7�w��A�ɧ��������:�Sg,��*(��d�����P���VQ.�{�@�H�:��'��'Z􀺅���m0�1����˜���u��gJnj{�7�i�j��+�ɍ"J<Yhѿ�)8U�gpH�:<�U�0�j5: n((�^q�?\��(�+�|v.�-U}�����6\��^b['{�%g>�Ѧ�s.gc��q��H�����00�:bO[��&���]����a�>�O����IE r�A�j���d�\m�y� W��6x��`TAo�2.��:�9bגa�R�6���Q����� �RѼ�zx�6,���,e�Xo�{�Q���D��������8�o��P��9��ÒUH72�Z:�Њ�Q_��k<$<�ܻ��ӣ����cQ`сm�er�+-�ќ���a#W����,�u�������<�I)�gQ�ǩlA�xxM��0&-!B�kK&��	�s�����v;|@��̨���%�Ⱥz;~X3��_�g܏ٿ&{���pUH�/<��*V6����Z}$MV\V���c�����`7=��Z�>�!@l����B��0Dk���o�f�a�$y���7Ȭ�-#����ñ#���x&�BJ�9p֔8(��l��|[�����r:�<�!v_���fYrN����Pc��b7��=\s�^	�ӄxa�/�s^�m�� ���A.���bٓ5��H\Nw����MC�0��Yd:���3ԥ:TJ�R����ڦ] ���k��1��L�5���j�[�(i��%*�<�5�[�����r��-U��x��_6at�"k�չ�=�:oH�"9� �x�[�x�t��8>�s��g�2�lR;?��:}��c�'�&�����ٸĥ}s�}�La��th6S��������Sr~�$�>0��0A�W�{��=j��k�Je�u�Q�Į�?0���Ji�&PR�����_�f�#z�=XlP�$���:�-=�?�����l�o���O�AV�ͳ֘`v?��y8&���ʀ�olə�]��&as������x�
��xl����m�~����L�����qPi՞~U�dyYWϪ��eS����Ǻ�d�T���9�Rqbϩ�p Qe@��ݎ�c���`&߄U ��� Ezote�Ö�������*�cE�n�������붮�Jļ�B�cq��\���J�;�.�̗)�N|&Tң�8@���74�oE^m7��-n���ڸ���L6`�!AD��Y� ��V���0���փd�MLX����-�M�Aw�ff��ԓ�4^}
�l2�Z�_W���}�H]�:p�!��w)�Uļkԋ]����Z2�G���)r)D��H,�!��߾<ߧ9u	�k�o{Qm(�"@m�&��Yv���y��6��"����i��r��3�g�k�Z˩������B��|`��2h���m&�u�K�৹��H[�^�l��W�)��H�+�K�ſs⧈���o�*,x4���7J��u�Ի�qW2`��0c��y���y�ْA��GWeJD��:>��l�U
U�Zk���[�ѫ����`��ʈ�c�^� KF�o�ր''wx�A�Y-��_��[ꁱ>������8��ހB�����=O�ãl59=��c�:?�S�$Z!D�ѻ�^F,Hy�71$)�U���5E�(�&W�y�+��:�3��jM���b�&H�
NM��J��%JE�,�-���:����J09�6�ci���k��"J���;$0�t�MԀkB~�}4���& }@�v������vw�@��E�I��$�f~썖\�<��g�d���������e���,�nS�v綣�����&P��v]��ș�8W��g�����.�}OVػ�1���2��E���_�x��� �Ê�C��W'1�U?� ʺ��J��RNw�|��G�����U�$b:��Y~l�-��4G]u�{����γ��>��jȕ%Cd��WRi� ��������\օO���u��˦�0��K��iY�Lo-���nV��߽�35q�z.g��`�o��0eNt(��v�`l�d�;n�e��˻�t�`+dS��*X߿��D���#LO��'���G�r�nY�z�dh��H�nU%�ј�ѝ�S`e���HT��le�iEnæ@+GO�E��i|Knσ;[j#ئ/T_��&b�2� ���R�q��N�AR��N��w��{��O%;����wnҏ�T���L����71�]��N�]^�:n��EA7�=�$��A����}c�m�J�<x�z��g��l��(�� e|�nFǈ�,�+�it���fLĄ�ð�ԧs�߱\���?u�@��P�d����R@�d5�g��(µ^�=i�F��ҥ`��7�e���Z�Z!���I��!�L����l�M�9+�<��#�}�(�	T��A��f<�RY��6��Q�-�)��njxd�<"ah>S|>�k���
��;�h�4�d2���/��.�MO-�^7�ҫ�&;	H�AD��JE����CT$�)����^Ѓ�R},�0"h��M)UN"� �(E��Th����:�)ƫ��y��/^[�u����i�W��D/�C���k�l�ޯ�
s�
0[��;<��-n�'���L�/�������^U��ͽ6�I	me�g���e��1U��{C�e�x�V��(�$�9y�Km��
�VƂ�%Ʋ��3ٙ���7l�`+�y	��5FZÎZC�sl��?p^����)��4*�.!�Cx�V�9�y�Ř���P�x�m.�n8�ߙЬYo����rmF�%�e�n���^���M��a�<|�m���7:BYQɭ�1��q��G��Uܳ�h\Q�?����uu����Û�ǁ������iˢ�W.�l�<@K�2��z0C@?e$�Jrm�S`2��\ޓ�䶳���g�(��9�B�;��N��@l�U�@�k�Ԙk�	�]O�}�xio}'.�������#	a�]zy�$����5�0�ڰ+OT7n��r��+�Im�W�!D/	�-�#��ؗ��回P$)-_'��4�s|���?��E��rrO�ʽ�{w����ә �/�3kN0?�U5��ޛO���Ph5��l�c2+c="lX)5@��XPֱ�`�a���a���w�i�y�%z��� `�!��ڏxuw�Z?�7U�\	�����H	�n�\U�XU�$�z�M�3p���G��!�m˻���CC1S�%3g��5h3k!�f^a��YZ����0V�V���\������D���׆^OfysA�;�o�~QR�s"�����{z�8*�!b����t_�l|⸘R����r�	KJ�D9��ae��3���������&{D*!|�G� ��͙����v��2�b�>�V�
��uB�_�>��S>X��&��y*��Jij��/e�NN}7�z�;����/���Ha'�
�^����f#��<Q��p\�X���o�6~�#�cY@ƍ���Ϯ�?�6��7
�@�",z��걪��o�φ��t+��%+�cp4���\S/Iu�Y?���L��j�X1�`�?�.4�>���̰�����[W�x�u?�)yAWUj��/Sx$<F�3ގ��_c|\8�#A�Y.�lp]afwSv��IM�������\�Ύ��)��,�F���
����L8�#副A�V�*������^����#unOt����߃e닣wI��:�#�Vh�I�ʀPӖ/m"�b�Z���9���8���w� �N��
�i������d*�c��^������Z����n��I1�}����ϥ����㦮�Q�yo���1h�nt��ު��<Hi/{�q�K-���+&���L�".{��r��A�{����{���Y�W�v�	h צ��a���9�����������`���!벚�/>�G����a&Z��-�`5�3�\�߅t����&{N�,�;qq���X"��c��o}�B.I%ɴ@�j�bs
2�6!ߣY%��?j/<���Ig,���Y�0�~��ɷ]�B*KU^$��Z*s9��"\��1STL[~��%y�uN2t��H���A�E�y�yߌOR<g�z�uq-��o�Ҥ%އd6�=XҖn@��49��4����/���l6�<�6:���ZO���$̲VXIPw�E��A��?7u��t(WT]�'U��t1��~�-[��u������L&���`�IP���H$H(߳�;z:�l��֑�_�.3��ӧ��8�Y��xX�6���X��ғ`��f𸇤�|��W���N���+)�~��B��h�^R�ЩqUw���s;g�?��'��յ�B��=N@�-�U��� ������u0O�` �0�L^�̙��[,yL9W�y�L��w�^�Zyi�@�¼Υ�uY��Fv�J?��Q���J�/�)m>��s��z�9INAF���E�5��*Fd��l/K����_ԓ\\�u��S0��S��\fy�>�	~����`�����)�0x$��YA��A�H�n8
ߩ��fk����ep�L��;iZ���-݃M]MyQ�M�Ĥ��K~���"IÖ�ǝ�A�)L�S/90��@��C8�����y~���-T��� ��]����6��t�xLs�!�]/�k2�IKN��q#�S.�o:�c
N[���Q��"׀͝�n�˔0Zxf*��[	����+�������ky�z���!Ϳ*�xj �Q*:l�����L9tlX��,��4�M9k&u����"a�����$�/���ՠ6� f�u��]#:Ɓ:�[!)�42�����H7, /�=W\7qC³PI���҄�-���1rУ�5ff>g���c���l�o �quO5ȭ�|�W���!�5y�]����0�l_൒�?k�5m�o�y��nNepы=T&�ʞݖ��-_�מ/	�ZH��n_uK��i�0�O�7�`��8�g�������D�z��ھ��,D��
}��Z�i� Y!���h�g���l30�)#tO\�x.]�Ełs�gљ�qUJ�
Y�O�[Rt��p�g�<ʫЪ/��5F��i΁%��{<��d��C����YQ�r}�w6����m�cf1&��Ί�A��h_�`sa6y�	�k�����-ߥ�RJ���'^�3J�C�Z5=� pKW��Ŷ�B��A��N֡��<<^��<&f�!gH���U�r�$���������R~�l�3��gO@�c)C��Ѓ��V`��y��E�|-E���?+��N��DQ#�H��-�$�{�Әc.,��s�魥V��P[�',DS[���9ix�R��c����7~h�h��D/g��I��� ��E���f����L�X����@����R����f4�Q[�	�P��3:yu��wf"��%����0/Q��R�}����b9���)̛S%���pi�~�xVL�Ҷ,b&m&�+g�w瓉֑��[��&ٌ�!�]V:�t���:&���"�<b+��B�5�($L��ε��"��Or�,7-��]��{�{��T��В(��or9Nk�H7R��e�A>���F��+:���NZ�.D�Q�22�>����g�\e(ڹ$]���IB;k�J�Z���ὴ19�4�li�T�.��j�й� ǉdE�;��������w�y�ԗ�~L�Н��kJ��c��Y��զLHT`�����|����Ӷc3ސ�*�	�s����3��0.T'.C������'�Vw�;n�u��'��r.{4�-*�݆$�§�Ơ�������T�G6��KF%4�Y��H	������=z�G�xf�-�-&qcD)Gvz0��9#0DkM���:.���N�' ��G�b��X=�a�Ɂ���X�n��-��y��$�$:�p�1�z����=ex!Q����+$f�����۞w�@�e&z.g���u�<���{=MQyi�x�(�'"�¾��=jjxkfؐwl2TƐ�`�@�b��wu�����_mJ�I �89�EGrW�Ql$����f�`r`�%��*jm��^��_8[��6� xM��1(L�u�Ca)��R>�.�>�d��Xʟ^�C��[g�!�|z������-S��X?�k�|���Ȝe��c�́�K��63����a�AN �윢��"���g��D�>� �C�.�?K���"W��Z8m�~�L;΅txP��d�G}��T'4:�o�1zbҹ�6�4<�Gfd�邸����z�z9��=c��4*4�}����]������-��rPu5�;�X�!'��Y���>ǵryS}�k-����:>>*�BnC�P��`L���H��\V�Հ���|������]�9�.�;�,��M���s��Q%ں���C�}֗>nj�HWJ�Vӧ�7��+ϋ�������h���^���%�ßV��6�k4S�ͤ�~H>�#��(Ϭ|�ݼUƜ��wd��A�m����`��^q���k}��J��{���8�wE��2��|�dΩ�axΌ
a9ǉ��#Y��R���m�D��I�.�Y\��p_�K����o��UtPa�:Q��4�"7H�eD��2Q5�f��KQ���'C���0$׉�����d-���,��]�ӈ��.XuV�f�Ìu�3㆜yr?��.H[������lPy����(�?,���� ���u}3���������Mrm�>*V��?L�����'��ِ�= hO�t�[�����DaثB�D
'$��&���c��'���_��{�!����"��yʼ3�n�+o{�!����U����k[��⓵�;Co��h%f��RF�-�Eڴ��74AW���5b�ʓ�!1���L�	 ����D�{N؅�#=+q)����D��+;V0�D�,^סA��El�+\��Ǯ�jxY�=�����ز��҃"s�`�jN�9$�r��ݹ�g�Vpi�m����Ś6.���c���O=Q'Mڂ�Ȕ5��4��Ι�dҀ��Cݢ�l5
�LWU���Z���frd2���[�B���V���=�)B)�N����@)T��;�U�CtJ�����h��aO��@�)t�?L����f�~�m�ᰆ:�ރ+��6g�</��6�d�� u��:�h��� ����S�Y���
�|�	k
�o+/wO���&d���>%9#��>@ъP��|��m]ͨ�h�̬��;h�B�L��.���i�/E���W��R�~85�j��:��R�R�A��^�$j��O`4�����%�z�J��3]��ak�R�6@ֿ[c��Rʫ�	
��(ꉆ]�a�y��p݁�WFZ��pBb���13e�Ǿq�O�A�oJ-^�و�|F�0�� Y�!�[���;{sl��tov �u���xC�hv�Xe�/^0���l����H�P�BMK<��M�\}k��8����%#W&���t��!	�Jdv�0P���U|����$u���cS>P�v!������� 	�;1vm���c��#�p�����jr�|��D���ɤ�l��`�S��u�'������	��1����P�����\4O�̩�1�;b�@��p@��x�۴K�c��&�4�fپ�=���BIe�� ���e)��l�(�r��MX���RB*]�+������X�^9le��6��)$
�m��0�"|������M>e�C��R��
ۚ��^&K��3#��j���0g��gPZŰ�Z������%����?J�ĭ���55����­c.\�}e�{�k��t��dJ(FL2��o�I���rI&�3q��\��`hH��e�t��n֫�3����X�p�7�9Ղ[U7k�S�h��A�L1b��&�"ǂ� "w]��"m�%7�Q����`%xM�e�C�I�Y ;��cy�C��H�~�w��R��x�U�]�@x��sN�h���+�P��`���s��e�_���ez�zD�����:�쿬+s��~�DoB�x7�&*��jw����E��8�J�c���'>z)36��]
�����}��3,1����&?>���Tv�]h�ۜi
�(J��j�fjx�:�����^�-�\�[�"�\��׭ErT� RI$W�VBg߲x�K��t���ӟnx�˻^︓j��h-�����׀G���A��|����I5Dv1d���7w�!3Wt؞ؒ�yy���'�=����p�B�̣��+`\�����Ҹ!�Ҩ�}k��H%��|��x����b�Xe�S��{�T�i�J������7�#諸����L�J���9_Z�F��n�$���Q���[��%��������4#J�n^� �+)ݿ
����.���-�I�kX�Z��;.���@��|ˉ����o�g?mW��Uw���?�y��V]v�,z��ה*�� ��	�mع4�K�����۷��!��̧�(��7��\�F��ZopP�)k�]���0͒`���^q��I�vRj�1��]N'�6 ����)�d����W�y��x�HLe 9�.�Eq����!�9�]ނ�ERѿ���\�!#��9
+��K��@u|�/�V꣘����:�vv]�$E�?�y�P��0��b
�`ɰ�ڑeoE��PA�K�8��`)�4n3*`�#<�{T='r�
���ya΄�B�����n����eB�����F)W5Mh�Ey/9�δ@��]	5��O�����S1 }���m˦�H����T����
���Р4(t.�Y&W�;�x��:��j�؛�[����-ͨ�p�h*�t��H�8�?���oK��ªR��|A����l�,JG ؒ�H^�'���o1��Q������h�,&D���%h	z��DHN�#	�~��.��)?B�d$��y��2F5z~V�q�h�@�u��+��\:�?����˃��;��������q��n��Re�$����E������*��$Y�6P#��ҍL��S��a@ek���P�5�������a�q�t��D�vo��d:�T8[�(� ��"�r�ڊ|cC�ќu(~�Lr�_C�����r�D̙M�79�j+wE54�8���"mj)�BD>r�)k���U~}�I_�ylg�u���U�s8���6�<J;�#��+h�fY��)�6�Ah����2��'7��QH4�`�����ȃʥ�B�RY�*��Ul�-b"�b\=K.���1I�Y%��vy�pԎOU�̠����K��� ���Ƶ���QȊ�����2p����ԋ��t���=	���a[��\�/�s,�"c��L����ߚ�T�xjg���\Li��y�c޿��"T ���P������v���A�͐��*s��J��^��7�C�C�O���2L�����^�Df�
��==s���׃/ �F.	�v0���\�ݳ�ڍy��@?����jc�U����R��yOSx ��4M�/I͸�R	��]���1��IB������Nצ���C��&��*o���M����(_��$mX_��8�fW��u�(��-u�JC���$�c׭�(����jF��/ \��u,�[+���[�mf�@��wT�:R?�
���o�W꾟+��b�Υq˔��0מ�}��7��� ϝ�2|�Ú���?J�ҋ�E��ӱ�(�E�ElE6�<#�Ҵj)�z����Z�Q���A`������%e���ty-]^l��X�A�|�b�}`���7<�1tI/��b��ΏZ�q .ޖª��*U: ?N�:_�����;�^F%$�w�ŎO�2��\}ם�&�s$V
y��@���ڂ?��c5*"�a��~��p[����ez��7�\��� �|�+���q�S��4\��n�Ή%A�=>u0�(Uq��<��~/�kl���s�2�R�Ǎ}�� ��
�/��&f
$��R�Q�^/�}ST�A2Iud@:�������WJ��vNH�0����i�6m���JN7�AI�K��ҿk���ڨ@�� p����_?}-����6��	�O��?�t�	���0�`|a�h��"e~����}D^Yet����������Ո�j�F;{��ٷWd�'���2�u���	�]ńh�ο�!?��T��C�A��fcoL�Ɣv�2�ހ��_s�6�L��sE�d�@*�KU��(L����⾔� C����������F�Rsrd�c�'�3#SpAq\{�v�k=����\�� i�@���'��{����n��$�Q�7�d���?1�Z��o�����b�Q�i#%�U�(.�[�=�#�����ST�AamXD�����s�����	B��l����w�bI^ݗ{SV�Xᒟ�EG(��Yp�9�4ǷR.Ŀc`N݊�1R̦q;f�E�ӎ*P�_#hH����]�0���;���B��ؕ�VAjᘙ���]��� E�\��ذs��C��F��_�eTU�\-
��k=H�QG����ɜ� <��,�ۇ�
'��؟c�g��:F/|�f��۪�%-��<�p�08�v"������� �ο}�YM�⣵���-���Lb�}N�ƻ�?F�s%�H"���*�M�m����p6/"�N$}߭����������UŬ��s�2��>�G�}h��VI�4ŵZ�xK�����
 :��'6���*w�����ƒ6��6��Z-x`���G��*PYA�<n^����wt��j�#��=��ry��U~AZ��!`�H�*�"�`�O��`�:+~³��u�w�'7F+\X�������ʦ��1hQ�b����T�e݊��g��Yi��q�07�U�p�L�N��J�u+I�Np�S�P�����x,�b�{���������Bԕ>5T&,ev�^O�9�V���!c�Mt�q$���c1x�fh�&�LV�%^��fX �8��O��o�v[x�w�=T�x[-���S2�fe�(\xl������OU$4�9�g�.S�h��qZ%�l�82����%�1�`�x�Z���M���L��z̚k�r��h�_r�<q���-���_�}��3����=����u
!b�]���C�Q`I�:5a���x�TȚ ����
?���֍�3��o�-��lj����!�W��nb�Z,2�'�rH����c=(+�G�c�w�5Mlp��sXA)��H V�p���^}Rk�U��&��6���i�W��c�l "�BZ-i��dYv��7�Υ�Ŗ�X������p����� �"�'U���5��g }ш��:/�:-��'̆�?=�?�N�c�;�!�����b`�9�c�j�wi�Cy:��U�ۑy7�q���_���(ξ>�����w�M���є��l��W��Ә�z�!��CՀeн\�}"�èK��HU� �?�o
����]�.X�#�\rd���j���ev�_.�g�����i�?O`Z>����w�����㻒�%�W:s�M�t�F��f��Jt�>ɭ�.�FA������>��t�x �&s�ډQ����mA8�u���x�7�Y6�=F���y���Wb�f��K�L��8�D����q�#�P�twf�8[��.�Oj�Νe�d�zD�����͞R��r5�R!�g������m��DFރ��{�q����xnl8��W�9��w������e��o�m�G��'�]/�[V�[R8���B�L"{�a$.Cbm1�DF?�q�C�U�s4�ĝE=��m�mUg'�zt耂~P�U]�����$5��A��Ҽ)�J�����@���q8,�ٰ�0�$&=`��훢
}w����甗1�>� ���*����YޤUV����5q�eaU���UE�I��<Ϟ��D��.�g�n�0����
|������t0���c���M����&����ՖC@�$���&l���m������[���=�P�1~��#��2{y{�Qɝ`���yyH�[�ez} &��C���{CW�F��x��F�rj���K��J�#�<+J!�v�F�W�$P{>�%0��Wa�U��^T�J�2Ef�Yͣ<|a����jf���^�}�c�����켌Y?y��a�~Z��c������/B��~C�C�|��i�g�B�Z�e�`�l�C+�� �t�#*˂jWE�Ru:�ܧ�t8n��
��e��>�Cc3�P=��� �����e�'3 ���t\��X�ʯ�G�N/�Aݾ�J�޴������N������{x�6���IJ�H��@̈����~�`�!��CP��qE��H��d��~㖎���2GŒ:&Ơ?������[�� �Ӄj����t,��dS��i��`��J��;�&g�j��
�9����m����Zߢ2���A�h�l�]��_S��w�m�*�ķNrd�Q��9KS˦B�� ��2���Y�\�ٮQ�0�}`e���P6�\C���l�&c�z�v���X�華I�+#;r�/�N��Ԓt��-�� Jl�PC�p�M��-��iż��\r\�X[���޼�v�E�;w;ZBu8�e����o��J���\H4��EU y)�}鲤�l*�sb����SƝ �D8��f6	��-��u��û3�n�+�1�Kl��>��&!Z8�0ɮ�A^,F<�E|�Lᯖ�1]�Pln:�N���#otn��5,��JK��-Adk��e��U*����GE_��&bS�Wz�0�e�����h>D{����~��@ʐl�}��&�#6�m��4�q����P�<j.^�*a,�@#o�i�A+K%��5�Iׯ	>�Z �K��=��j�G��i�_��\Oy݊u�c����gH������7���kN����^cv4`΍�J�V�uӦ�<�%<|Qm�}���eGZ�-l�gw������7�ӊV�$�����&!���s2��w�zV���Vi��Q׭�7�Y����q�I����~'� �@w�<��l��q�����i��!��\����}d����{�5�բ驤�yqw�as�
}�M]��F&]N�����4/�������I^�L����x�%�7,|͖�6�q��9��mYeLA�A�8�	�+��`�����p����"�����_A�e�P�)R��.������R	��ඊ����M9�}��7sm�&���a�n�B*}6��{d\��# ����-|��ӝ;c�Ä�]�#��zh�zCPs�k�)��ﯓO����T�(��=�V�O+�w�Sb�dy8�׮GP�{C�W�/h8�ML�#)|{��n��oúL�bZ\`��3��|t���)�� ��^k�@׎"�q��!<K�ɪ'bnr96*��KӞ��ڢ��2]���'��:���~aX`�׼º%|��\-�/�w����vU�f�$:C�)̼d]B����	����C�J����Q�kV�E�%p�vhm9�"so|��# ���+�'����}ӝ�Z](�Z%�eC ���9��95&�M�DK:����~�X�~�!�%=1��N�A����3%NةxzB�T��q}�W��Z-��Cƹ��!j:�3�i���F	e,K����F��ꛨ�{s��=��r����cg� ���7�u4��#o��� c� ���X4iݱB U�xF���߇��<L@7 �uc` V�jV3�n�.�Z���(�Ҏ),.I�ߍT�5/�
�٘�� �3g)7��G��ҋiw�˦�5ܜ����)J�4"����*��ZZ�=t/ѳ�����>�H�JS��������o�Ù7����
��@R���;!;��i���w�Q6���##��^���abh�.�Ȋ�<���S���� �@: ����)�����Ɇ�b�ÿzi$��3]�"�/!�3�yHm��
����x�d��a#Fd:����u�|�F���/���uf��º��vD}ˢǹUj��¹p���x�Ja:^�Q�e�|��N�«�`�+���F��y��u���z�[g�](�^\�����)��7���сM#Zg�fc0����������Z���ڌ����U���� �>b�r�e���tߣ@M�K��|W�E�͜��;��E�?h#����N����a諩;X���y.G�p;��Ud���ǻ׋�����W�Kws����X��M��{:e���|�@T�,)c4�����k-�H�y�D
����Dw��5��� ���[�@�z�a���IH#����k@b)�@��-K��a���	�M/�����x]cV�JΨh���,�hf�|0uʰǐ��g�p�8��E"�W>�H�ۻ��z�"U��<�'��h�!��D��B��bZQ[������D��R�W ��<df{� +f��ε�z ��$[EtB�\�9�Y��? vw������Se�SR8�?�C��������W(�`�n��:r��+�j,ԅ���l�G{�8��n����O�
�^��6{�|���k��J0O�x���T,���Ճr�+�r�1�g����,s[�:p���~$C�j0��R�0����~�I�yp���d����wc����0�&�~Tk�k��6�q�{��m����{I��P,xH��	���Wd���X8��4����'�g:{��j�iئ� 
��*vl��5�C׻G0�<���x(V��C~�.��Y����;�^X'@4��W_;>��_o�N���H#��VdkZ`̩)i��S��{�C�X�Z��k�z�V���uu�(T�]�8s�����YA��HyEry"l+�YM��߶�J��a�i��V�bQ��, o�DO�L�~p� �H��rȡF��s��zOv.���ܷ�! ��r��dO�d�]\�Hc~([o�W ��/{vpcƉ�v����A��b���1NJ�$^�>頯�z|�4mH3��:v.�n�/�v�j�e�m�|�.�`������N�%'�/4�DGL'{�����!���TSA�U*V�Y2#O���'�uVN� i�ZRaյ��R�(
#Ŧ�I�.�(4��� ﹈?`#d������	�Q�3���!�ƻ�?��F������*����MK���I�
��,��]{��c�%(�ɭ�s�zH�����z�nmgDM�H�H�m���� �4��;���5v�zN���8�$��A���n1�"�f,_�~?:�E1]N�g3��_9/�Ɲ�x�Xh:����;�p�]:5o��Hѣ1�7|9V���G�Ds��u�������`���7Piq�빠�$Ded-�C\z>�b����`aȷx7��=�cM�.$!o��c7�H|"1n^�i8)��ˎA5��t����0��e-�	��0wU�*�Y�f�n����y���a\����`z�o��\70Z/�zJ�f���V؞�@�dG-2�O��T��`�ro%�xN�-_R����J�W�:��6�����)̲l��
g�'2�2��3�� o���J��ä�$�N� ��0�ס��r�,|��~�ےg���y�"f�,���x�?����!�NL���r��
D,�x��[ӯ⍑�e��N7��)�t)t���ׯ�����[E�R��I�����nU�S��?'W�Es���qN��';[��UKq�ّ�=}9����K���+��qM �u�7���͟�z ��l�Z�6g�f�� �+n�a5�.����S�Wi�2�^C��0�fUqp@{���.�c>�z�d���!��,~�[Q�l��ju����Fr��������F��Y�#Ȅ��g�I��cNynSr����]!�30pE�Y~��^�kfKփ����y\�:����Z���nyCr|DxM�֠�^�?e��;����H@	�AM"�L5e]k3T��(s���.�U=l����
2t�]�p�������o�~%�z���iZn@���l��]����(�D$�n"��ʰ��αgʵ���7M��	��C���$y�u 	dv	���b��q\���7?��o�:�=����PE�I�ϼ ��s�,lj"���V����~��qC�G�����4'�Ȧ^�5��!Hx��C<���x
��kj�]�r9�I�*@}{:_0\�-��I�<�6��U�BA>z���1�������p����#ޣ+OL�W�;>�b��Y"��G����ɉ��i���&'F����� cL~�%�ߗ`.]N�ea�"*�䐄�3�ҽ�m`����E�������.ȆCQ�5�Z	��|ɢ�2vC}H�5�`� ����TE�>�,,�;�����6�jY�E�`���OD%N?�	J~ڎ�_n��so�H�`��_�0�C��
�
5#�U?=Z��Z$D�����{쎴�gl�3�Hu�5\�$�()6���%����v؇J:�M������/�ա��9�<ŋeC.%���[;�o��7ϩt�^-��D1��f��Ō3� эo����X`�G�aG�$1V�����
_�2c�D�֮��o-�?w���^����	��v*o��85J4`�%���q�n�f'�2�����A���!�Ъ5��'כPS�nf�o9'1y�r-%Y��e��.��ޙM�[CL*�i�E��G;k"�?���m������T���� [����XBő-.��A��T喭֏~+��q
����%�!y��.���׽�B^��۩��{���xNݺ�`3��.�(#8	��+�5��ZC#��.ˀ����0��'��7���ـ�����Z���L�rH�
P�k��� 	aeY�����=����3��t�l�Ձ�=|�Y,Rū�+���W�'�4��Sܵ���/�R	s��'��|FC��ޏ��߯���=�i�Z�����/#���{W����Ӫ�L&Z�- �)�5zÜ��R�% �U1�M���cAt��B���ws��6�v�&u�Y���� cHP��# G>�nF5v>	9��[�%.	�J��Z����c|�?^a<N����
2��"EQ�.@�1�>ȗ����s�~����@�ԎO�5 �RXwa��E�=\�%���@"ӧ�1Ch��j�&��@䟪�d'-�1n�5���������#sQw}��qv^��0�U�R�¦,��?v��j�<?o
�m\�T�$ܙ�ҁ4�7�A�p����C���u��pl�����:W�X�����ҙ�;أJ���F��#�w$���M��Qf�,i1\�f4�}�6b/�ɧ�Y�S�������u+�1e�՜q�]
�q
��p�D�����:#T5��:���?W@���C��<8�u�-2{ַ�����������G�<-ZnY�:�*GVg�>׺v;��ny�b���J25,����A�r�n�E6��A��7�����N�c��jc���o��\������5��>�'��2��-����b��a�N���"���,W�i��!޵�\���
Mb}4��"Y$&�-�T�NՇ���8�WU��J|�\W+A�trmv�8��""d�8.z��� ����	Iz�UvT�� G�_a �,��R�kW�g(��dq��1%|�� ���k�O�;�U+�LJ�2&�� )&�&Rѱ��D���>���E�1@�@��u�+�J�>���:���rW@%��e��NN>��.��,����� )���}���A���H>B����T�$�5O@��2�:gb�C�	�x��%�|�71�sONf��^�+�L�o�0r�_ڛ�֖`)2���fIm�!E����K�a=8E]hB� g�o@nH�x�U?l��T2;����Q�V	~'<����������f9�Wb�KV�. �x@��g���|�Bdf���A�k�-�N��3m"Y����޺�&t�1��x=ӒQ-7:����Q���P�gY6�lv���}���'�2|S�0�̋�bP�z������q�ৼ�44�j'��F<�F��4 D�����&������w���o���pB����0Ц-Qq�����/� ����k�9_�ksڢԎ{�xxţ��`Y�ž���}.��Br,�-v�D��0û��G���_n{���G?pļ`lџ���|�9e�rٔ{��-L}b4u�(s7��{Ex���s�>E;���L�T�x���&>w�[N/1������V�0�\�}\�pg
kA �]��-Z����Q�W�"������$=���-4��XbG�m�$"ϕ�ڢƐ��^��l@�#*-����5X%�������j�^)��L'�P���������:�lQ[k�P^�S���P1Ej�V1B�d�k��,����>��Tcc�xT���-�qU�zx�D�C_�]H���05�ֿQd<��}~��S�3JD�#���"l8lXv��@��[WI�R�r��bA��KUj�@7�Q#<�^e� L�;'�^p	Y3�	�5�$j���i���$����9�Vp��G�K4ۛAN![��[�e�������NW�[���=N�ķ��k22�t�����Z�A����Aj\GP����^,@��v�;M-ݟ��1p�Fԁܭ�)��S����P]��i����	�#�^R,���<��
�NH��D$SB���	��7��힡D
2`м��t�! �L�7�ju�G]��e��RO��T����4�
&67��?��ME�!*���.����@�{h_/:���y
�N6����[�_��S�fbѰ����zz���x�9Y��d����|�����N�"���'P�+��ŭ�ף�9~؃��u��/�jd��@j\�s\?A�.YfJ�&�]gO2������μ�'}~��^F�#[f��孈�� ��f5c2��JQ�̰���s`�<���냷�K$��@I��_efz]c#rLP��ԕ�\%�luGM�*��D�ۚ���������� m�V�܎�I�I4J}��2dN����p�/%,����;2~ ��H�#������N4��x�A3.��fp$?�������k�2�㮀_����5rR�K`�o,v��8�jH�d�Ȗ	bNe(���"RN I�R5�e�Z�s������M{�61���Ȉ������~qY�`b�o�mh#;_D)�޿�����.���<���;eC�;2ū�ɍ _�z�ns�Q�f<i��[
2g?�&��PpD����OEe��܂��D'`gb������t�Ձ�v��5��;Pe�u����donW7��R�{�Z
�3��1���ǯuR�N�:�ٱ�$���N���z��[~�~�e����ڹ��������9��	<CdO����Md�����=�J���#�뼃mǺlw�F�t�|�푲:D�
��W��d b���/{N厥1�/}c)��NAlHF��A�=�4��]�&S�_:Ҏr�:lR���u�5�"\߁�NͦЌ�{5�R��*A@2=k_+�9��ג�=��A�=տt����/�� -���q��y��`v�x�X؄}:`�%�>��F˖�"u���>$��.J� `��lTME����#�I1��Yr�o"�N&��ϑ�U��p_,dB���F�"��:����G�L�=RK<}6�#q��pI�m;�Đ-m�84����j�x��h_�����⑉b<dz���f��T����5��I��@��H*C�1l���$��=Z��9K�������e(w�:^��J�z�˥�7w�Z+�[�����_A�#e�N����Q�����g_H)u�c���>��>/��Ѧ�50����+"���p��5W������t�e"/Q|��� ��&�|����BB�~ge���]�	�w�T�@C�B��6.�W�<�h`�#׿�/"k��-O�M�g�[e'c���`�=B��=��bq�:x���Ȯ
>C���֑||͚3��ElY�b��ӗ�ų�W�������W<�(�����%Q�/)��7���･!xP=�|I��SD�qO�1q�N��Na�b�m�pr�'ώ�>�����X�S��B	+�'HoP��|V�g3n�[�i�����6�2�|/>*�Q��<S�ԃ������ɤ�_���B�Uز����7��^蒦��G�Q��a�O(<߫r��1�D�e��L�k��D��Ո��M��˅7�N��٨{	��V��5�MrY7��֏,e��q $��>��|������c�^Ҙ|���N�c6-�B�*Y��>���A�+F� �G��ma��VE�n2c�w������D'��JY�[~.�4��M~qMבI'���a �sq����>�����m��<}c�/9�(D��PK��wt���k���Mf�^����q�'s��-���uK���s6QB��z�i�C��2� �UՇ
w��������4T���~��o�	�̵�,�rp?���G�	��
��YR+��Y������wP`��6v���i���EMU��,�A�_aW��w� �8M5���Ft'@|���H����&���i��#"\��j��$��;���P,ڜ���6����-�dRp��!8�~���Ɋ��J3��%�Of�Vgac#�/�&�Ԁ(��M�~�Ei�7�<�Cp�{`ե�P{a�7�p5�`@�`^W��/�z�A�jC�H�qb��W���C�-���OT���(�42��z��W:^�nT��0��O��ֈ<�뙕��m���~��ѯ�9�U��=�f�G����q�T�7�e��/�|���B8���X��&Z��]nk�-B�4�g�&
4H���Z���M��E���]H]tA|I݂S���,�����@�M�~��%��1%,�jN�O��Wy�F$��Š��bV��L����q���jB�.aNo�l�i5��kFE�N N���A'�m���[�Q�G�B���2�զv趸�o�m��Nvm�����D��f�:�@��:^?Ơ/�V�n���PIE��%\E���u�Ot-��{<�HVC\V��-�y��*�W5�_<�GV����_������VR��@FL���#�I�f����\�pR�c���F��kg�0ҰM����G��e��P�Wg��E,G�#	)�6{d(3��0��b�y�l{7�	4�́��C��M������׈�V�h�?�Jm��*{��n];U�XEx�k[�G[�Lb20IY�}��h]�ˑ�QS�����c������� ��B��Q΋���p��e��x]7���Xo�e�6aflj< Yh^��8�&M�w��TQ"A�lF�����,��!�d��|B2�Amv�+ML�����~���4I���6��7Np�FYƂd�ST�����?7���)}�%콁��"�Z�Q`a�|Xe�����_�!�4�v�V���V��އ�3������c.��b�(��%۫���D�r?)�@.�cxx�,�7-��Np�O#�N�G�m���L�޷����sU�@����v�@N���J���zя�+M���r���ϰxP%Q��!��E� �թRz���Iqn�f�}>]���t�H�����L΂'U�y�E X�4+/3����jR���7LQ�?����5���:;ȝ�8��=���6�u�6��ځĚR�qYǨQB,�%}Š�K<:r�QM�PB*#����n��&`���bf	V��4b��m��_�\|�({:T馑�iSъW�j��g
?B�2��}S�y��Api���.I&�2���H �?+z�d̑�}G66�:8e ��X�GKD�ډ�?ђ������.����a���"M	ʩO*��1��zS�>�߾�T����m�)��������r�@j��k>�*e�W5Z<��>`Q��}B�8P� ���d8��q.L�ҼD�=	[���ŕ����jt���-໌F4�c��_@.u$�,7�X��bp���a������e�9��w�;��Ó�dO9�<,)X��N[��I��t��\<4� �G:e�5�x�-��ØI�_QC���,PH�iy���P�'��cp��Gc}y[��S���J�?> V��{e�R��o^�/��w��iW�F���L;9����W�q�*�->x$��hI*0��3p�%sy���gcٞn2�����$��ev�Wnj�"9<�1^�+
�ME�G����D�����@W���)//
���]�j�ù��6x:�uK�/�Xx�q�:��D�;���Vy�,�j�����І:�/�8�����yD���{B?����uM9����}��Y߿:�%�� �Ku���7��{G)"A8�����p[_H��h��i��>�K�����zM;?\�n���p��>�v���3���$]X��s�`��S�+�����w�Mf�v'#���d̓	�_u�B) �0����2O2�9ԫ����Pq�Ǝɏ��'T�W	�].%:�B�%��I�<i7M0�\j�W%��ȫ�L��(���%g�|�!���JG�>�yt}JckAٽT���Ȇ!��eA��g�^��RCZ3��k��l<=���K-����Iy�Á��(�/�����#�Qc��H(�l{�͏
�-���tf�\I04#�MA8��/M �����u$$-�N�e�.���l�jy�p�]�UaM<���Kc M̀��+p����n���v�n�� �t>_ �#ق�_�o?yOqЃe�������� �l2�2d�������ےe�~���ޞ#9�AV(�2p,{Af�_��ȅ�v� ��g��c�*9�n�9�}�4��s	�䛃�?qx���_��[��K�6z��:n/ݟi�=�D������ ث{�v���u�>`�\��b.�oi�U(���Ye�d�?e���p��g���*�Dm�1ܬ��N���N��Z��y�fe%3UN�]�Ha�Q�s��6=R"v�I�C([HP'B��4k�R�2�˗y;�MV1��ߒ����"���,��;�˓~!�6eeR�`sJ{&�{������JejQ��ؠ&�bt���l��ϒ<�й����&���#��4���H�y�,A��"�K��:�K�W��>D�l��r��v�o ��� �y�n�2L7"u���J�Ǵt��a�,
b�gS6��U�Nr23�~�C2���"=���-f����{V����S��a�?�e|��sT����� �y�b�$,vg��f"�ԏ9��[j� �ـ��]���q�;��d�6۶�uGz|�U��K"��{�]�O�Gl���/��.$]�Y�e{x���\{`T���X�̇��-
�����S�U�V����=�	Ѯ��T�|��T�!A��
��lY�����%q��%�~;�m�V:.r�\�{$Tq7��e�ʟ�\��
�������sk�^��#���Z�-g�2���p9�<�J{����}���l��;��2)쥄�a~)Z�a�[Ws���X-��QS��HW]��U9Ɓ�J��J!&)HM��3a�bs^�������|} 9��6�e
iȁ��tk;������ŷ �=�
��
���ɬj�Qz\m����4q�����7�'g3T=<��Y�\�ig8H0'SS�_�b�ԡT]�ni���4�Vl�B`��{���A���������i��b��^�B&�Ր���N����������D�v}��y)o����_xbPm;�c7��5�'֧��1��{��=���*X�z!���pҔ,�5N���}Ƨ��ŶlF~���K���Q8'1&+�~֦�e#�
��M����+�F{2m8��݆g4pQҥJ��bз[Fb��񏗼3X��sk����bf=\��9��vLI9�q�(����,�~'��F/vq��L���r�<Ճ�3|j�S���E��A�?�j�H׉���|��`?��=)[F0Ex�e%�O�� mwN����ͯ�T��]-���N�#�B��iʃ9��.#�!Dz֥���WƓ���Sf�w�f�A��H����с�Mԣ�����.J	 �R� ��T!=���!#�����`��Ӊe�JE��ů�R�_�Fx�*0��8r|n�yB�tw4ÊCVR���l���d��%��Q@���Z�Z�(O3-�Q4Q��m?�H�?���p:���o��q?9��2E^e�;1<�i(����S���ӈY�D��ɑ}���S���ns����\TfL�D��޺���~��8<�L��9�7!|vo�rX��A��9�;�҆��cԽ���Ϳ�3^�(��̥ň����J��c`�'��f��~XL��2��7�Z��}_�gW�y�?{'W?`]�x�e.H�5�Hظľ���y$%ދ��`���kR1�Q������Jf J�y��ϓ_�H��2z�EQ2k����8�,���f�������ޠx'"&Fpp��+5�&�<��w�UB`���\��I�̆�%@���.{��Y�{����NV��վ>�A���m?ޛD�[Ld�Ey���(w����D�Y�Kǳs�D^>
�O��m���R��������3Y^�*�*CO�R݈�*fl#��*�a���0��?����67���yLeyk�Ǌ��נJ9�e�~�h�/���l��ư���n�o�&!�B0�u(a2Rb�IIpS��&�8F���'}L��߹5S.t���i=��M_��<�OU_Y.,K*��0��.�v�؜[�t��\�����`/r��Fz��]tt{/���x]�W�¥�A��}����ֈ9���ҋF�⛶h���&��v�{��\�o��n֏��)ڑ*���i�^<�9�X��zi��n���w���[�4H����+�Q��e��LF�����N�bY3V��hhY=|]-�Wd��[�}h2�X1�rܒ�=�M���{�\���i-���b��Xz`��zc�3�����A)*a���xHJ��U�V�����o�����UWaY-���3����F��a;j�~���}�~!'pͫa�36��w�yf5np�\�wv\`Yx�6$�lG�N��JQ��%���,���3tk���4@78?e��s՜P���o;��@d���@E�KF����~z��~)��s���N�	�f%�� DR(,� (]�����lˬ��\z�����~�JQl�����w2�ㅡ�ER}~O{+������^}���,'�ӆ�T����0��=���STr��ׂ��\K_��#�v�������4�^�`�H�L�v	�1����P���n��
�wzm��1 a����"�3i�g�a���Ճ7����`&IU�%V�:�l��UC�d"���( ��=�y��\��*tÓ�kW0�pє_����"_Q��$��H!y@��gW�4�w���I�&B�ܒOp_ �Jmm��h�|R�KIH4S	R�L�+��uf���9~�E�4���%$y�Z����=b�˛!F�1���{�����U��FР��ukDhdnm��t�����ṍLv��4 ��Cc���Ё�����!O�`X�}�i��&9y?[��ø��!^Z�t������������>[��Uī��E/�mq����D3�օ�Ξ:�����pJj|O&V��c�:�7��6��{�oڪ3����_/�����Yz�}�7���۴  �YC筕����rޓ���!���u���W!u}/k3�d+�W�$.Z(�]2Z;2k$ߍY�
��%(e��ɰ!��4.��2���YOH����9���
�u�b�+B�'&�  _K�
��C�1a��C�cU��ʛ%�@���l8��|��a>���57�d�F�n��(a&�5�*�d�0��>x<_ݶ���pwGM�n����;����ǂūv�q����w/ĞG�D�cc��Ŕ��r���*5��8���	�����1���Y��ٮ�!)NH�[l/c¬�?�/z��g;���P�ԅ�܊$\
#8�W8�lX�Y|�yYS���-��}�i)$\�,X��W��f���גe�?�XY�y?�K�_ug��KF��t�C[��=^e=v�p����_I	��?���!L��E'�Ϭh0�U%Ә�«&��5�a�F��E79}n�Aň�MN�*{��rȈ�zf0�tj�[i�M�h�5�p�nLT�{yq�� A�'ni�
&z�?�s��K�~�g���R(���}r!��@9b���2�c��ifEb^�6ٗ�R#i�_�i��I�Z�框{��(o�౅G�d�6i�2�cIl����.�w�̑`���4�{;�sl�5��n���}�֬'�8>�7�e����������a�a��/F�S��ٻ�5T���.S�Z�7�zO�"���#�Cj�0��ι��WP�L�O���PyOd�J��Ǎ��+�A�������9f���> �$�el��v�F��$���=.l�?��b61�Y����X@�P���F�u��Dʥ��=����a�<m��,y�藑L�B��Ed�G&�騏S	�NpI},� *����˞�M-�j2Lx��o�W�a��@���js��%�ץ-�-�D.�V�F�-;$JpY�t������b�b6'��֣�t֔hYj]�D�!)�ǒ�^uC����.>Իs��;��"��>s�}�p��iDg���0�;��S3+���k��lj�h$�RD��1�����J��tP!�5n�
��/���%�E��/��Ӆ]V�[;[ (Ƒ��xS1T_��Wt�b�����0π�o���n�4�W@�����1q�̎|�f��Ǫ�Z[�e�!�y�۩=��L+�uHhb�^�r����Es�K[�7F��J>ɔ��JP�;���6/���O�cT��U�誨��zX�1���}/R�r��P���EǏ0[��P{̼6��}�Y�qf�jI���v4M�eP��AY��+�s��[S����9kQ~�S��A]�,�W��4�φ᎜uSXh�a@��>nebTZ�Uw�*+�U�3M��Պ��ӌK~٣T"����YSTO5����^����MJU$X U#Es�v���9�_T~�G��t���"�Ɔ��qGr�H`V��u���k��a���qE`2�f�t1Ԃf}�5��K�̌4��Y�Ț�*������@�]>�#���5Л����V�� Չ@��O�&�QG��9C���(�ܐ���骃4Ѓz�d��Swg��<=ŕ�����u!!��r�04l{�aC>b�O��#B��j�[K��6ߣN7F�.'$����m;��0��<������U
�[���Zm\J��Tc��d3d�w�j�blݰ�R{��,*����CУ�')ćbJ�i?���pPC_
�B��ɞ������f<����p������G�d۔fO21!�kk���#��ǿ��\�7����`D��Rr����j]�*��=e�Y���K� fmcS���]���[E��v�G/��:me�@�%WX�i_���6���ΨIip ����B|��EN�u)���5^�؆��q�#b"�v���{����V}���diAJ��ߦ����Qi����??�w�[I݅��$ui�,#\}���,�>��l�\�@��h%�~�!B�-���(���f	ٺ�O����A��>��c�q`О8�6+��ݙ�����`�CQ��������s �0ځS8_{[��@��Cu~b�z�������+��p�KH��������s�T�����/!� N7`�f��K/�T���щᕉ�w��/�D�T!���7W�ѵ�/�� ,��	���,^ �;���+���/�uqм˥'��6�u;�y����݊l�K~�"�.^�ly�0v� ��&���UM*��ϊ#�	y��H[4\�z�Ɍ7�>���Q���mNX��<H�Zړu��fX+�͊D�F��<�߲N ���kZ�%fb�IJ|�ؑ<��;�ͼ���H���9��<�V�e�ԅTT����0o=���bn976��Pg9C�ye����A���(ؙ��OU�?��b�I������q�
�I�0�t�I�?T����FY]l��BK`Kq!Iڮ@�k���a4��E7��1q����z!�u�a�(�eƞ�E�&�O���FQ��M���Z�ʚKA�xY�@k0�v��ɩp�^^w
�E������oP�c%�<ǯ�:�:4'�P%����z��ݶ	�I~}%�G�l,p���' ���t�[�_T��V�i�`$j�ڜ���ljM�I,���(,� =xt8v�k��>'�ѮD�����˰P��3~E���0�U�4�O8�`���;ٴ�U�_��.J|�y56��Q�¢(��G��ٕ�5�"Hrfz�>ÿ3|��R\�}�a6�7�D� ņjA����U��{�9��տ�"q�\�� ��C�w��g�4G��A���#��?nqm�������5"�%J}����"�E�9��~����RWƓ>0j7��7Q�� �[���� [VD�;���2`�-��5uH���TTm)���c�}z�a�V�CPA�jF��w |����o�ᕢ���c����# �ޟ �@#.��*��c�2�|�{�-��M6 ?��SS�+�?z���=����o;:� �~�g�SQµ��RoA@����M���� +J�*���nMi���e0C+]^��6s��3PQ�F��=32S?���K[s��^���?c�e㯴�T�6zp3����W^7a�
�^C���#��:��
�?����Azբ	�f��>ß�%���S��Q�.}?Mwd ��Ĝ��3TP�,	K�I��k֋{���H�AR߯�d�
��4L��ǔ���LD,��:�3�T�!f�c�������Պ�ϭx���B��Bh�u���U ����)2+�X|����~s�,o��ä��Ga���qz��=���n�I鵌��|�G��G��J�(ة�7�C�F���P�{�>�RPU"ߎZ�~w�� �$���м�B��^�l���9�p���E o�^W��s� �@�M��qv�Һ#j��v0���gw0Ԑ�hZ���R��CF�c6�4l켋K
���O�u��]/���i�^��n��J��lO����o�t��X��hQk}9�۰Ͽ�R�S�.s��3�����p�:��iq��n��\¬� ��g���ηwyi�\	�-�TntV��	z��ϔ�GnH�Y�����@ ���`c�K�wuuz�.�:�9�� �*�]�(]p4K�O�������q���K�h�В�!8��dP'�����Aꊓ������V��^�{����\OlD�揔^���V;]�E��`�B{ �-2���'B>�(j&�Ӎ[�(J/��g��C�/!g���vs��r�DF_��x�4puZ��)2H�͒����-�?��g*������I5Qc�o��vs�	���e� �͋r��&RF)��w�;���$�d��u�3[re��z���wC թ	O�7��9VH�]$��G�o9S���v��G�)�-gw|�=,����0�ت�ͼ���J���¸�-Q�O�N�d�!��u蜀��)ml�J�S
_��
��c9VF�*"���17n������w�Dvo+�JWW�.q�A���lId:��s2��>M6� -ja��\5\�D ������h�|��� ����BC�C���zpV��(m��lk��t�La����5�@��}$& �����e��a�����2G\��Eh��0�dv�)��ܕQ����$�z_��\�W?��(���k�mI�:6m�d�9!-�/(�z��E�Mވ��� ��4Ӟ�E02*�hP�����Y���i��I��>Q��Z ��P\*���S݅�\�m��CV�ݠ��}�o��µ^'5�V�	#J�7�7�筶��܇j_��VQd���@��){J�T�[4%<2A��4�g�w�=�X�ܥ����®��NC�'�U��mD���,��ҙF܎3'��̋ʖL��1�V���_h�yxa��˘x��ϻ���?_��U�G���L��CI"@��L���%�̐և�_*�_���ȴ���Di�3�ñЂ`I���/��>�qCOV��/�l)���
�u�>O�P��<z�)06�o��@Y,�k�(*=hԘ��U������uD�[j4��,D���:�c(�\�����Q�`���T}E$���`�qP��*T�VR�V:��bG�2z�U�]w��y:q���T��?
#FigF��>:��Es�(\�4R���θ^Dz�P��G�h\6�Ҕ �� ��!�H�����D�2�%�vҞ]�`ʺ��t��H�s���^�ɳ�Ӗ�U�ΰQ^ !���%��Vc�x���7���n>l�=\�Ga�k��QE��'��I,�G��
Y���@lHV��S�Ć�G�/�S���ڙa�+z0���BSi{9@�`?��"��#[�'�ơS�󉯀h�JzzCsה��/�ݤ%'4�=͐'��32.9q������"|�4uʀ8#g�x:6<t�V�w��'
X�mhl�ڧQ�P7�E��Μ�SU��gh�[w�����B�s�͓
���f/
{���uۥ�;M8�7��Ύ3��&&!�YkF��}Zd���\#���|��rg�:X�&���ꆆi���"=�ɍD=���ܱu�>�#�;��\K���_�B	k]֩3+7M�EQK?���//���V n4ER��	'�h=��+��M�i��2� �ş�]Q��AYp�|ý�f(�]�Ս~��!y�6Տ�>���j���r��}�Oq?�L(���O�\�A�kK�3�A��a� �,��Mk��6�~�pF c�.�%)$ɣ1��T!gԽ��8�v#��鱽Y�k�=��Pg��Ir }t&4n�˧k����J
�`d8��"�K6�$�s������2�q�-ao֓��(�x��8���#t��.��e��*R�HS��H��^�;��N�JǸy�F`{�j}qˌ�f=�2��#�h!!7nSp�8�)�_�lƙ��Q� ?���3704w�f�9��u��b����lX���@*�zN�L��l[�ꅘ���| m�o��@y��d���e
?�+�t ��&�v:��O2��R�#I�0�R*z\�.Y�6v/��c'��$� O�D�������hK����ֿ︩�V�3F	``еR��8;|��pYҽɭ�rpr!ZA�w���7t���@8`B����<|iB5/�ɤ����QO�=O��?�;���	�Ժ.wN|���6N�"_K�b���e��ӗ%|�!�<@�.8#�p�����c����jT�/<���#{����d��/�ϻT��E7��y}�yţ�֚ZN�Ix�i�E�{؝��D�sŕ�D\��U�Hg��&��OZ�>�R��=�R:z��T��;��n��cˮ�\�fK
k�$�9��Q�#8^�Xw��2���MՋl�+YCL,�/���ss[��+cW�SH���[UWeOH�C���9|l�Ɵ���>rَ�m�#��:1�3�O�`0)�@����Ʃٍ�����g�$���L����x�HU(��B�}�
��_A���l#�����ᡶ�"�z��1����W�?�7 �Z}�=)��a����}'�=�˩K.����J�5ka�B��Cĸ��5{�5��}TcK*%�~�^ �젊z���w�Cn��2Pm$
]�(�m�d�'�	A�����?0�=���һ?^� q�0�[s/��Hyp!%Ф8��;>R�	��Ytݚ"ކ� �t8	�..�kq>�$%R�ҷI~�F�=�&|�s�,V�
H��-��$+���ԌΏh����<z�\��l��/RTR�;��]HK��Q,����<W,ǘ��Om�;LPf쑯��}��'�+S�r&A�4>A�"�(E�#�G����:�;hp�Ng�C~m��K��4ԇh��Mz�I�7��[�L(:�J����
�  �������pZ>��.�����-C-(5��C/�Q���qN���}g�Q@�2-�Ӣ_�7�U��x$���M\���5-=
�v�%Cec����kо�Dv�i��2ִQ���m�Y�Hl?����Z��3�8�,8�����(iؕ��l�o]�-�d&W��e���г�'�F�>�3�R���+�*�G��Gz1�����q�דo�3W�NR�Y�'s-�󓖒<����挙���/�Ёú��B���瀔���!+ �  ���ڋ�hҰ�Z'_��W����<)��O�vȸ�x�r�9�GQ�%GU��P�њBJc�����x}��-�eU�qa�Cc�
$�LC)[�H

"�<�~09�1�������{�h�_�����(�g/�(���]I'bX�7�b0�	��7$�o������,^���X��i�~�łR�!pH`W��6���M�l�"0�)�:uGA�$�
�V˔�+��h�	�Ri�%� [gIu5���w�B�1p�#W�n�#2��M���ut��&���J�l����_E�z8��V�Xg�`w���4��Z�������#�P6S�΃UhU�u�dq�MZ;&L��C,e�/�G(��#�L�JK��~vsݜ�u�*���lr�5��JǨ�{�S�@@�B[u�t5N-kkB�/'��Tg�C�G_ľlgK��WU��(7f�?�����y���S̨1�L�HTD'�K����\��`���캗�}Qᯇ�v�W0)v�ğ�#��bA�_H'R�g�:"���b���d�3�&����I�,�Ci�P]����tX�W���ݔ����T�Z~%�.a~�9��e�N(���m��n�X�Sě����ƨ9ܲ���`
3�9y~I Jd�$B�S��-��pE�mu	T��(�}ަ�IQYH�lْ�9io�1#����gU�8����(+ׯ���E�g���e���K޶����d聚��6�Ί*߯��dl�ꇑ*�ܟR�D��`e-��:{ڬy�nj�KT�뒆Ǔ�����*N��nn�7�ۓ"Ȱi2S�п���<��-��;>�hԉ���ޟNn�e�8���g�x cfT�>��l�W���-.�mhm�bv���Ժ�_�N�
"C�$Q+�$��'�,D�Y>�T���� �j#+b�Gj)�
���mga��<3�N��R�\g��4�LЂx&��k��%�� �-.e��peAt�K㇫�t/�Y�1� N����%i��O��v����v�9�x����[��yk��!:7��/p_5���
{�Z�,ff�C�w�r�rm��3�f��Cǂ�6��O佡e����d�"��AUM��ݞn��;���.�ڎ���b��Z����/�8^�5�x53�n`�J}��&�+��;J�x�<��;R�nڑ�h���k){޾٫��6O�s�� �^�����u<�\B����e�A]�G�q\81P~�`BY�Q��p5��A5�?�Mv_��q��"{m�D���=i�N����ŦuC��:,�[ba�	��#���9�T;pa�J����ۇe��i�ޢu����I������Q�(��f'�&N�}�;�H�{R�J=
^���s�Cf��v��`�H
�ݮc�O�ܢ4�GFS��"�7���s���b����j��kVNbq�U�	����ۢ^�p��1�(����`)��<���;��)&NUaTy��8?��)�Lx�8l���P::F�f�<�O¥�J���G�b&Q����\w5{�ӹ���d`�-��	p��?G���c�z0ٹ�����A����@M+ �ϙ889��ES{���/!�ފa��Z)�d]W�*<"]�,��>'�v���31A�т&����lSh��̔���'Ǣ��(_\�5
��#ttBw��S㠼����`J��~��tL�k�rI��zŜ���T��4z��c}���wْ^Q���Ŀ?�X�b\z�e�0	����M��mKd�Ko`AX"M��:���A�L�P[3$��t��ʴe[��"ϖP|)}�JS���9!��}��͎ąe�SN���F�t|7�de���5�^�~��(2&�9�Q����gg���W� �5�9�[Kt���9n?3'�֥����ߋ��3�'Ů}[k�wU&Cb`^[$]+��<����݂�E�Y
���x\?
Z����u��{F�]�9�����w����79�b������Ooi�	��h_���I�[ޕ�7���u����kQ|(p��TS�H'Y]K�V�?����8��0�h)�J����ݘ�g���˼�
ce=>t9��Zޙ4#}r��03���=z�����؄��P��rٓV)��E}Z�$�Z�B��5�GT<��NԄ:�i<�h�4���r�ܐWo�M��ܫ=�]VB� ���bLp���tj�m;R�U|3Es��M5X���q]fOg))���Pf��i!y�.FBUGBv�~ȥyP�6$B��>[���s����.����_���?��k������߹�Xz�ѵ
����a�l�a#�9��jt��I�w5�)������.��e��>� "x�G�ٹR�U%Sц���K�*8w�應�k�%��Z8�C|��Z\l�~���ԏ���
��D�-�.��^�fj�^���_pw`�'0Y! ����g�)�n���Յ]��&�T\�GS�8�������/� :�qL�"ZQ�<W? �ȍ�?Ľu��<��,Rנ���<�Y�j|6�0��J&�[KX�ro2+ilL��4'F7?;��@Pب��4�eDCP�$��&1���6d�P����ہΙvӕ}l�k;���4��Y�i�e�'�O��r�"�TB� Z�y���(�u�&ؚMo�z�~�o�Ϸ��S֧lS@��g�p�D8��l�+��@��D9;��z`��Ɍ�Q�>�̤᪰r���X\�6�#�HFǯ�r�L�$o#S�L����y�p���]�u���0��`�]�@����+}u9�@C����{�H/���Ui�������War}ĿnZF��_��8�+g�[*5�.,�*�{�g�r�#�*&&i!;nx�F�#s�,gh�j�b��7ѝ���H��	����[�c!�5z��u2�����E�O
e��p2��B0���A铊w���P�Q���E���<�H��	e�������g������D��E��5�/�F��FF^3�-&�S��c���RR��1���\��,=R�6������rNT�ҋ�'0[�
���"~����0�ms�T4$��N��hb(��iOCo���b��)�`���m��~��<".a��'L{V���a�K�>� "U���Ӄ�,����"Cu)̟��]6hs��pc���������T���@�^���w�,�7{.SfYr9�����H�Oh��/�n��ڠ_5�0�GVj�D�CnQ_p��
4&��bj�>U�T��d��Mj�L,��?�S�z�
%U��ŦWE�yRP���bٗ��L�Г�����Ȯk�=З�ÝL=X���kQ^_�Y��ܗ��&�^���͊V��_I�8�Ћ�"<{ G�uO�<�6�a�%�|-�k�k�.ªO�VX7E�<�~�T��)�'�ǈ�P�����~	��C� 3/�r>#�;w����
6-����;��s�<ԅ�7���x����k_��Jx�zT~�[�=�O9Ǌ�%��)�ԻY��w��D��F$�s)>�((����O���@��Q���W
����VbH��^���6 :�5P߳#�;1�{2����/)Z�f��?��ADUpB�8�Ӟ^��}� nN7���p�ds��&Њ4��a�c������v�͈����nb���s�c
$Q"��r%�ռNg�~�B��� �~�t�;t�Q��X��q�E1��A|��}�`��}O '��̔'	|�n*�hIu���i���iuE�Q	��9��Y�ʗW���!��gMp��R~m	�ڴ�_�[�V����I�qC1�Gpڔ2��b��	Bɽ���*���"��MNd�+�,i�ho;�*ծ!�p}�1��*�Mr�]DjmE%�|m�`#�,A��l}�*ξ�Iqc*6���1��w�]ty&�����w ����W��!+��� ��]��]����E� �!�1�{��ԫ&�%(k3d�,H�r��E��������t5�˼�S%�_q;+��v�Ѭ��7�M������|�p�L),�_:�T����vНY���T7X���Z�L-�s�-K�����%t�i��#zc���c�-6��C���p�޻, G\z�vt=� / 3l�-�c�^i�?���OpSżK
�J�F�|�P�֊��6>@=���-�]}_Ƞ	�x�� <�!�����S�ȍJ�q�'��K�	���CO���������$����������6��(d�W�)aE1Ml��LI�z��9U̬�7P�(Ys�S\M92�I�l@�S��fD�K,��b�'����'{�k�'�XS-��ЖU��d3�ܱ .��>��I�ԝw̞�ga.H�d��w<y!T͍���$�g` 3O��bB��z �?+��M����e�W�5��;��[�L�[��k��;u�9Q����?#ۏ�	*�7>
�g�Ⱟ-��������>�D�	!4��P��@S�-o�m���5�HP��(�9���i���w%ъ�O:ry�H�f���g(�V[!�Z	������F0��S�1����ӫ�)�qP}������v	A�Z��*�닑���W�����f����ZK�bUr��O	��G_���Hړֹ_sRT��ԕ�/�,oq���5�^u�p�L�=p�y����κF��^�
��&���P[l���t$Ң{G ���8�4�a�^�E{��s7)c`K��A�*H�X���o���#pQ
��������I�/l�54�C+
w�ӨS̍���K�% ɱ��ä~"�����,\�߮�xW����p�u�\;Y�	=ީw�7�#}���9���p��I ^h�D�ޚ�,C>̐���V��lwM��S�pF�N~190s�<Y�v.��Rm�
�f�I��j7��?@&���\1��;_�Ӓӿw�����`�Dur�}oO�ө�����y��7�����s�L1��q� �w�״�H;m�<�C�u����G�\��)�����C�s5-�NHX
"IˉE\�?	��ꊌ�8v����CDF����E�����x�ׁ���t.d-kP0+����Zw.�x�o�`أRRT|�B�6��@r��yF���Z��rXڡI��
�t��N`H
���{�(k$���z����S ��z��r�"f�޿|���E+�zʼ#�9C��"���)C�Fj�Wh�88�w0[����l�N�9�6���L@Y���֙l��}C�?�k�ڥ��~EX<r��i���CE"+��ר�a��r�Rm���`�~��mʽ2�b^��,P93#�"4�=x`�zGqsc՟x��_js
���h����W��D)V�4z��В���0aOyf?>��+�ޭU��wR@E���/�[��Y)��O�Cn���瘫��*��)|��r���"�V3�*i�����r0��y�K�)��6�)n��U`�Ez���'���tue�K��sVL���_V���V�{�z1ٻ;a�rSg(#�M��\���^ï�W��ﮜ���)�:Ⴭ�z~�{���-1�5� o���PA�<u`�g��=\ǧ�hW/
���y(����E��m�U��PL��K�}��U��W��{@uU�W�o�1���(����4�[�XK5�b%�M6���$2������:�3hZ�d����T��ʩ1���Bi�˲��/��T�	�ُ�Z��OةV���	:�{�aB�M��u7����SA���{��V�#����Пv˙��4Ɋ�f�\���53?�i�'.�,�7f��`�P8��k(����U���J�_>�!�"��j��^��Ig6���|�Ǵ��h��V���(s�v�4� *��?(
�/���~�t
d|$N��9�3virjn��ro�������0�"�)����V!Efn��>+�~AkÆ�W�P�AA�^�o���~���lFk�s=�j�؟�n��L����"{69_�mZn�VR2��s � ���pe���_78��iLԢ��UM��Ʌ�g�	��P�2)� ���/�b�.�)q�� L�V��D �z�f�����MI5_�q�u�y�ɹ?C�dU�.A
��e�"��s��7a�(�ʜ���X����b)��l�'�3���~E���D��DH���!23�Bf�hC��S�d�v3J�&�ˍ��d�'��=���g�X��D[|���*��x��JpH�8�Kb8��dj����JCqlnTS�{�;�	��W.N�CmFZO�7Q���}��4ߥ/}I�@�"Ə��V/Kk�=1�ᚖ���NƯ6��IZK�f��{�>���7�@$��򱹮kig�C����ٗM���.�s�I
���1϶H��4,/pIXs�i)b������x��۽�ו�=��t]�Z�˴��x�J��1gn�GU ��\b�e���3@�ԻK����ϓ?�Osm����_.��!x���+���6�	><e��� d\�@ƙS�Iԅa6ٌ�e@��c�=����k�&b�P?��
)~�}�� �6��Z�2�M��JY�a�X�+}e�$4lz2?dmy(�]R�l�������v�=�D��jo�X�=�4:Q7!��K ��E���:�3ϻ�[v=�/��qbqD.�~ �v�����F3s�����H?u��* ��u����(->�y��_Z� x��[���s���%D��,������7(����0�fC��l �t-S����>Ub��)�u����0�5�9��;nQEE�ؘ�O��<�¥�S�:1J�M���d�p̊9A�*좝��A\�$�CxP�09���T#��zʭX^j���:���#�-@&� fa8,il�5���-�����n���lӞyDF/��i+�ɬ���!I���T^|�e�u�d�k�E���f��i�����/Kk�]�_���/�|�F��\6A1�8�y^�1�u�|˨Ɗ���gqE���[/@���<
��XG4$��Ft���\�d,uh_��L�x�0�Ij�'���w~����tD�gv@�h�u�Ĕ�;ؔ��=W���J�O��ѷ�GzK��bK6�U3L�s��E��o<N@�i��\ݸ+���Z?lc������c��O������lO�rĉ�n�B[}%+���0GY�Lδ® �������}���@��tQ�t1��Tm�þ������p5�yO����ml�&w>��x�ΖNC�LRH3M����f3؀x���؇% ��4W�㤐�i���d���ň��F�Ѩ*����r��tI%~�: �]Um�UL��{����c̓O�8���r͗r��WG�����hr��:Q�.����$8�D�}Zڇ��Kڠ�����Y���:G�0&J:%�>!�����v7b�wt����ba���6P}۩th���q\!K]�<����u��:&�xOk9�ѩ]P�Jq�|"��������?6�[)2 �3���8rO�|~:�$���?�D�y�lslgk��	q7H�K�"MC���3B���ɀ��^���g�pvd^�9�ڷR�x�C6+6��  3�+,. ���d7�o��� O���T�M��l%SI�/D���;��+��)�b����h��jl��@�_��3�LIq�v��z�����%��@��T�~l�����R?��B���Pt-�؁GId�C�/��$j�-ZX������z��͢���9y��:K?����K�!ʱ��_T܃@i2�t֯Uq�/mۀ�{"����
��o��%2��F:7u�,�g�~@�|�q�Fz����������g�=Np|x�1!ҝ$p��Kآ��h6�C�'��&�v�Y�/�1�����P�.WP"O�1u#�� Z_���j ���$D� �m��aO�0���-I�V��)+���ao��$~��_��e�L`����k�|l.ؗInGC����+C�\��5ҖIY\삅
���#j#%�q.FS��[�� �g�|�㷼��͂���J>GK���1,��+�Z�i���-6Ka�jkG�/X[_?m�\1eW[��˰bK�m��E�./����I�|i�x#�.��bvﱙEŧ��/D�F�h�]�����;P�l!u'��b�/�5�g���"��o_�����~��u��Y�y��<B��*�;��0�'
�4�28nj�*3R�fP戒�S����Ne\BWpچ�ۈ�2qv��n�����m�+��_,J�o��U��8JT>���˛�^�[>!�����-$�c��~hN�d�t��Za��Q��޻�6�'n�׳��Uefפ��$=��f����:����nFœ���lܠ��\����:k�=$�2�Z(�%��@���q �/a�<A���ֆ��b񅌙K�5m�JTÖ�`!��KE��*�zXHy� 3"	 �vip(P�u� ^�l����L��A��b��p���hb�KJ8�Ԙ`:��K�ď����H>�F\(���F7��LQ�F���  �5Ә�$V�߹'z�wV����r�J�#He8t�j���J ���ɻ�lw�ui�e��#UBnA����T�9��	�%�٣N[��m�i����כCv��(�ntV��/���z]f���/؋���j�9^�3^H.�	���CD��������;���ˈx]��Uoڸ�m��>�3�	0K��}F\�
T���������V��AO��H=�V�N� �BK�a?._������^�o3���F��?�=�벒B����a0+����mB��S`H���Q�t¶�i� K
A"5�w$ |�Z�}	��� �,@>�;�y���������a�%�C��λ�'�h|&A
?"�Ɛy#7���se9�i�Tp�~�s'A�M��$��T�vڛ^Q�hY�5˰��d��ώ���]�EUs�w�e��Z��9쓴�uT>���ʞ��6U���S��Va[t�hK���NJ)5��I������o����x��������M�[�P����f� �����Ʌ�[�k�������z���M�N���yhE��a��Lg�<�E�v�C�L�h�k�>�����ӊ=��:�E~��]���'�������{o��ً���~6*nY8������,Y�0+ŝ.���ƪ��ޗ��AXҶų?��ڻ�H�P��z4�� �(����qř��H��x��ژͷ�0!�+)@Q(&9 �HR���ɪ��R1�K4�.���x��-0��B"�ny�_:ϯ6j�q׺I�4��V���L��qT���Y���7���Ǡ���hT�p����ۇ0�5[X:6A��
˹Ca�Bu�� ����#��U��U{hK�wy.�4J�јPdLA�C�&h���ڥ`HQ!��1�*��=���i�U~���w���X�n9�O{��5A�.��j*|���;�5��<>|�\aĢ�"��dU�M*A�7��vES�_����լX���ޓ�������n����`���	����� �#+'�|U����R���)��o�Vƃ_�%*�S7H��x���D΃�������2xaU@�
t�}��kH��_�E�c�a�e�j��Rq3�g�A��Эc����4����(��.r$��õ7�΀4�w�/Vub뚍�z�c�����r�~
��Z��
�������%�ϢC�gg^�"cu�s RDv͏�_�_m��|X.��3�s\��(��wU^��!��,f�%U�{�OP��uY�RB�ԋ�2��	?��w�s
�k�.�L�6��_Oj�ď/��	8��|��~�c��e������c���1n�)�
�Y5"���h�YZ�L���g�������*T��C!���1�_��p쵸�&)��0/�RP��0�G��G�O��^I>�9���;^Ǐ��9y�e���9a�+"��Dlc�P�	7�^:���p���K�����+���'ݴF��9��x��p
��(f��x���p)���%+{;n��y��R_�.q�hĢ��6M�M�}d���s��Sp1�Bv��wa�ϛ5��()�F��
E�!9Cy��3�/#��h".���YnX޲v>�mߞS<�܉�V��>#�Tz��e����p�20 93q͵څ�(�J�tb�
��z��e�C���)�j��v�|��{m�k�V�a�Q[�Պ�Mkq~�+��t$��c�?Z���}��<e��]E�ty�9j�fT~3���8�/X7��#����֓sһ�ݣx�5���D=����
;�vMM:*u[mHw/q�CWUq�c&�9UOE�@����7���P�_x;�H�c��8��axЮ��V�Uv�^-�@����LO�!����s\`�T6BlK��}�9jF���8�K��P��ɡQ�䒹�9��佱)�bፋ�����/�X���G���%��ƨ����k[���!���^l��w�n����6���3��:�:�d�Տ�ݸ�w9�ـ�m5�H�"6;d���Y��E\$h_����Z�DNT3w��s�5��(9�6R*F	�=�,&�ODd���ƜjY��9�]���|��|�����X���״;mW"�+mq�~J���m�԰S�o��3.����9�������TQI�a��T��I5@��v�	��-m0�'3:KQ�m(Nq~��3�'m���
�!�u�k?o��z�B��	'_9z�[���vt����0�"������;������*�N���v�	���P��y����l�(�w�h���d��d����d�I��cz{��U�ƣ��W�����?Σ+� P��Ŏ��q�qH�PfX��'��gOX��Z��cQ̵�{�F���;Y3��pM<�>G��}4�W����	nwTdJJ4͆��ҺZX����U��|u�8e_���A�}xPqoeW.O�ID�7�9"�V�Ȧ���%&^C�����}39o�Ft���I��C<�C�d��*�v e���ЗA�l��sdB3K�5 ��>.��I��7k�� Y͈N:��<$s�q@�BX)hBRJ�_]N�
*�RޫH����&����T�^��kwGϺ�d^���c���+��E�I��U��5I}���t>�zbX�1TO�)Y�e�jV��W���d��2�N�D`'�6-���Q�>�����X�o(��4�����Q�@ѣ���u&�=Bj��^խ�!��o�al������m�_���o����A(	�̵�ITz-�`	��T�1m�f$��yK-��,�(���,ij�oPB1<_0��F-�<��[���q&�d@�}j�>�°���-��$��£�X<1�%�ʤ�hN�	�Q�|W�D12�Dt��M�T�w�ca�J�å�h���M8J�:O}e�D�`��{"Q����,NB�z\��M��$�U��'��B|,gIW(�1È���P�f��N[���x�Q��9|��"d�(#\����L��k��f��?���ͽ�6��\����
u\��’vに�9�qҽ7�L�`ޮ`zR,C�����k}���H�A����w7�ĉ��q���1Ob:S��1𐶨R����ּ����&#��v�������ԙ!�'����f�W%꣚#�sʽ�O�T� �"�mv�c���aC92������B)�Cv�Q��-<,�i�#g3#����Yw�,XZ9H����������jPi6�?}e�=��9����pNt6Z�S5�_�����\�E���Ѱ9�A�B�|0�ME[�}e�\5͎OB�?��K��)���u�T�P���vSO�i��Ӵ;,�[m
����\�ڔ�t���*�����aw�f�[�/���(��MT�5ʌL�O��`34^:Ɲ��h�T�]#�4�4����)��<����V	������ʩ��w"�`�.�:piw�4�W.�z0�}6A[X6��^��1D�~a���x��2�z�g�I:���	�e�؛�^��L�M���f8oum�f��p8����=�-_�GX�V[WK�-΃��`m��C&N�iN�۰�����7�doUև2��M|S�εd��jR.\J�cx:n=�꼹2?��ݿ���[L;�q�;�x��͈+��"X�#�^��V���B6|�����
�T^E�Ć@�_xL�'u��P��[B1[��LT���_%� �n���_�<�_�;��2I�h�kx�a���YSъ"�A���|�xH
��q=��&2=�{5`�� ?�7t�}�I}	�&+��pݡM��,��O8t�wq�A��I6��/uYeV�m�b���g5��ۖ&Ud\����>�*ݓ@
3��Q#�-^�^���_�W������*��7�%g��@!AZ�ħ\Z�9���I'tl���kh?�D%���]>g�	��mf!������P����z����1{�>j�r%�D�`<w����������ح���#����-�dM)�������]�߶:�o�wX�}�C`����r����c�Xsl�������U���l
	~����9*Ơ��xJ7n�u:5w5+x<�
���3���I~3B���3����V1�����Z	a�гX�A�]7��yZܪ��q��C?���mЃE�u�2����i�Hȑ#���W��.���m�Ͼc(�	&V�&�+�n�A�!� ��w@c��b�:Y�C���[�N��X�
�M�~#�f($˫��K�M���"Ond��e�+Y��{)��Y}H%FZk��3��ƾ��̣�q��5o�H�0��B1���̅���{ó��QwL��#�$v�a��� V��E��?����wt���_@�md���F����dyh�	�@r*8іr,�&F��#w*W�cq�J�G.|��q���@�2�F�D���Q�0������8%h��
O�_���� P�L�?lp�֚�I)�?��C�Q�v�^A��T���D�<rB��I�"~p,�)��hZY ��t^�=�]v�hgX���Jٟ�ͳ�qڦ��[�i6��`�����"��l�b�A]���]޷����!���t��<M��;*b0�����Z���=������J���S)Yrs����"��}J�Yza�E7��a�� �{-�:�6x�g�[�����9�o��-�W���5�D�W`U��1#e����_! L}�hwnX�ݶ���gR�z,RF��\��1J6IY6bk%�e��W�v�n��T�D�&N��m�t���0~���b�*;�A	}�{�Q@�C���������,���Z�=/zRH���!jx�n1�M�����d�$T�v-����}�Kj�)d����]��/.�WY 3������GEp��No-����z�ϥ
y=�̈��u����-V�V�/�D��"�ʲ�O/`�?㖭��V��1]Bq�Zj��<�bi���|I�1N>1�	)��SO.��W����_��:�;�d�5~�zO8�d,Hnl�&!�A7|`�y(Qi���n'*��{�.6��>��?�6��>�*�o����ws
��;^
��w��%��҂�p��n�r��璏���0U�;�#=Zb�ҳ���.���lVb�����
x�^�]G�)�e7F��lo�T��⿿HC��ί�k��0Qf��f�:b�g�;�G1�֥ߚ��;/�e�l�i�OS�1�($P^��)q}���'3T������6�b@�׼�G�or�ҟۅ�86�5s������� ��.���{oݥ�
c"�{߯n����g�]6�K�d�#��(%��"�d��y���;��D�1G6\�z%/N_���;{��=̯����/����4������� Y�hk8�ꥏ���T?�a��a����2p_������&f9��T�b���K|�?��U�ս����].�ľ|�?�/K��ĔG@�ô~�0x)�i��G�V�D{N569�F�A��TbVI;c�]�P��m�I(��l@+ض�/#n�M;F�Md�o�X�3J�?�}���01\\�rXW�GHx�V �L��|��}��i�*nNb�=��g������Y�
c��qZ�Z��3�" �ǫ�����[�*�TڛX ,�k���m��a�HS%U��=�'/uv±F������SAP��G{
I�'�;j��L�^�JZd1��_���;|� @\�M{�5����S���Q=/��B�#�);6�!dH��~��#Ҭv�Du\e����U[�T�rP&}UKm�����u����.���n��Ə����)��=<�C'�\eTbg���dg^��H�,��f%�BRU}���p:vdD�9����! �mx�2s-pe�.�|��!�ZB�xHX��m�F߬4W�d�r�6R���U��;W��)Wdh/��צ�Y����;�p���JS7϶ev.7�m'D�M�K�n��Z���{������>��t���ޟ���{ i=I��:��a���XO�ar�9/���%�	��]�͏��yN	�� �D�w"<��x:�V�4yޛQ0IC���#`r�a�
f�"�/��DF����am�X4�#�ìQ�8nݤ&!������d�5��H��ĢL52 ��\�k��� k���l�4��R���me�հW��Nu�Ϯ�U�>SΏ_Ѫ�T�xS�{���a�1���^�r5/���:��u����	�Q���s���͊��n��G`q-Q�J��{I��K�K�ζ��qJTjh�8�[nG��RU��yC�IE�ʫ�����e�h��U{5πG�Ҷ1 ��Z�{)��KN�{�|y������?���R e�NH�º����ޡ�ޡ��<O�g]����%�d����)�6����������0��E�A�W���U�_Τ&��a��Rk��z�7�^*1 +ܪ�gP�Y�Dۧ�������uʡ�HE�CF�L���������k{�!��u)�䐛U�;_�Iޡ2��1���i#��fY��$�����=?��j��n��*Ĕ�NmN�2op)ү��i���w�K��I�:↘_1�pI�NѦ�OU"�8�V�*�4ϱ:�1g�f���P�����a�j��*���9Ҝ�g�Y�s����
��b�D���i��g7�����r20Qj	Jbi�#s�H����e���l3u���mmǪ4	�_H�{�7,|�
v�.��X,�S}�c[?�B-nўҲ��Ξ)�pX�s���LZrt�����҇yثA��j���9�ۧ]�y���6�q�oc��d]�|��*ܖ�1�[8�'���P�z	5��ά���Y�(��W�8��6�Ioh���cB�����Lu��[	rt�`lpG�&JleE�˟�`Rc�E����g���D��O�����F<�gP=+�Bǥ�:��ײ��<���BB�[a�I���
��պ�:��h����$�4���~�Y��E]-��̌^M��L�����}i]��
+����\۞n9 �[��1�Zbv��.��ZXbW�`��0���^'��R��F�w�d�dU3f���q��P+?�\����Ң��iʕ���T��2�O���TXGܡ���3t�?���Rb="���Yg$�(���[a���~&�4���b�&x���V�6*h�%��?���T�r�'I�n�K//�9I���L˱�~Z��7�wSFosz�"�;d���+F�uYbt_�BvԄ��������b�R��8-k2�����j�5�T��}�����1s�����Hm�dV(�.�@����T����� 0mw�C7�i����kx����k��2D?��XH�"���z�Er˓�Θ����j�,���d��S��/b�U�:��Ma�T�ۈy��C��"����n��$�<�=HJڮ�vz �I�Q�@8��1�:�&�Q��+b�Z�K��9%ZĹ�n��Z/��)�;�G�*j���q��P�r�= R�]F�aUY�F��d!Z8T�'�ēC}*�I�� ~��U�L'yk�kX��&�1?���M��1eO�l��t��cF�7OI#�9��)g-�CY�ܢ�G4ν�G2ZBԫ��5��IM��*���)EF�q]C�0��������j�͒�5�,ї�C#�`� n���gպM,q�Wi����O&ۅRI�\A�߷%	^<q��m��ϛ���wh�9�8}q�X���T�q�:V�	a{R\���\$���(���R��0����R��߃�%�BҚ��p�S$�I�j�A|�ɭ�bY��'	��J��$��~c`	�*S��F٤ַ��^ug����P�U�9����zZ�O`�ݟ��lAk����=�A�p7��nF$bTq���]��n�F�dr��j�<ط������߆����������lS-;� Q��V��{��#W�4S�G�r���+�.<�1�$�ɞ��*ẻ�l+�aU�PȖ��x����N0��]%7�!�4s���dQ[���̈Ѳ!tZ\���G8ڃ��a�y�9���8����6m��y�9M���R}E��;j�;��$T����l���r���%��}=�_�/iBi9�갍��)3Q��(]��}�N��DE�U�5�lK�R����H�J�]t��_��x�ǋ X�>4� 2�mB�+�Kƌ�Օ�:�U���2�l�`K�q  D�Z2�NJta��B9����ў3�^*�w�_�b����-� �9��u���:x�(AI�D��q�J�y�6���$(dp���u~��u���S��
��A��n����?iͦ�P�]�(d��N��`i��d�Y������7���4m��a�O�Wب�!�KZh^]�(A+���G���윷�����L���+�4�Ԡ�G�P�_�J-����΃�0:�İd	��j�^=Kހ�F���� fO�����KY��J����W��^�ȁW�3�8�����F:����T�L��A���HA����W?��H�ƌ�'l�9���x5�W抛�;���߁��t�@Lj!�݆�a�0�+9!q�v*����G�j-;#�Z�vÄ;^ �̸�L7o��"��Yh��]�>����?a�y'b�4��fB������6 zz4���Y2�V��h��������" �i��
�=�W|��Zj	���(��9;%����{L���h��r��ad'��V�,y��ϛ.�E������-��.-W\���*�r�ɶ䢏�洯��[���#�'೎eaKޠN��dƈ����ws��x��(���Ji��\>�w^���|��ؒfJ5��3��E���&&/��SC���<M�K��څ�bZN�ڄ�{+��HS��/ ���'��b�-�́�8�&�qe���y�����Q��щ�F�\�S_�bb���� Y��Ҋ�G��6��P�{�X�pdo顠Pѡ�P�UN՟E�'�W�`H��^jf|���s���Mw2խ�M���S�m�'_Γ�*z*s����|���"z��$J$iЭ��؀���2�5�,����ǝ2�oWJ콒�$�U��i�j�����nᲒG�9��e/P�풧<}8��ob�]�9˲S\�� �y�r7JXd_=c���^��8��&kX-|3e�^!1����`�(
�&�����B�K��G��'[���#�1�Y�I1��g���)�F�H��6�#~�Q���˚�ݧ�d������~y9>�m�G�dq���'�p��v���A�PH6C���Y�ߖ���z�҇��(����F_0�9+ik��b�ӽ�,d2Ο7A�<te(S�YX�I�V�ӄ����$�S�XY��0m�hGV�e�dbqyD��a����C�4��ߦa�	�UW6���O�Q�J�<�1*�c���\#h��j�CX#��s�:��0_:��ȁ�ΔY��-h|\�"�Eϥʌ�\���ܧ�0���ia�=;y-���P\ɚ�vW��ѫ�b�a��J�����W�d��/��A�3��)H�apI�����w) �舅�;=�%*wcB�o}�s�w w�q�fE�
�f�(k^I���is��o	`s��M@���P �8�#8u �i�SY����_�ŵQ���ӯ���
�X��������X�f�T?%l�8C��n'�3x)���u�^p�E�u����.�7@�L����&�?��F,4~QV������}'���=��!1t��v���N�n!��������g��A�)C�� [��v\R|��5���$���ǁ01YٖR��6\�����ذ��%ne������BǢ؄�vq�����U�3Zp�ɱ�0�*����z���2�F��Yĝ�lG�	1��,n��ztF�$t�??�AU�e�mK�k�Vg?�4���t���C����h_�����n^S���+����jc��5c�q��5� �F�#�;�I\�3�m�=��b�~��<d{��_��I���7�B���1Rt�Y��!�)���?Ϛ/�"���~�#kġ���>�iA���� E��Xp<iiO��)��=8)hn�j�����4Lbе ��iYD�´w�FYD��h�y�SK�%�q���Ε��r�G�����Nb�w�_u�zh�Iw����ή����FLv�x��B�3��uҰ9N����Eɂ��'�^�ދnrn�8����i/3���N�]QBk�⍰����&�H�Z�k�3s�+7S��۰��y�P+LZgpNj����$������V<9�l����%����a�����+����c��ݿ[���]Z�e~�A9E�K�ō��(�~�)���%�Y�Y�(^��*��.3����(H�o�S$}C��;;�7�����h��K�:�v��e;D�xJ��&lS�։j�i>/�=��M{"r�	����nY��(q�ۇ���uj�3pu��y�����p+��ݽ�z� j��̚!��)˵9A����3r~���h��N8��7�c�><���[�.���ih�1��X޺��^G�)/�L)�c]�%E�J�`z�]�p��9�+����,�����7���CQ�a�~^3H�V��;��u�(�5� d*#T+��?�Qzħ�0<����7�H�?�uVn�b:D[,�����s�~/���.
���S�wӓG
�`]Zg�YO��H��)�_���4w��N���j�����4�[6ps_��ŕ4�O/A,�����C�j���e�:�H��� `��k#�ĭo���\G�G��	  0ˈg)6�*ջ�?� L�w�'����SJ@Kd�<t����z/F9��7�WR��]�xR\e)���Z+bGT�j�oGHe���P��iM?�<����"���,`g[��[�s ���35���3�+s����i��043Zʷ4�m|;�ۑ�����y:���e�w�j��ץ��I��S*��: Z1�ܪ�����ܣ���h�.��'n*�e��Z.�����G�R$�c����`��^������t���)�_��?8L5���	���MRo����^֚^w�X-�M���wa���ɥ�z�ܘx٩�:�A��T}�p;��֟�G�9�Gy�n�!��W9���S}Ag�'O1�b���(*�E"�є�(t ]P������[f)�����ŀ(�ע^O��F��m�Q�[N"�Rd���_��`eA��H���	rpZ���pQ�t�W��k�I�=M���w��`��Q��e��k�lu��F�,�=�◢�m�����T�T:��DuP�4�
�OX�Bh2��"�������녫��Wh�lt�`�(b�4@�^��C��$��ZEN��hgޓTju4ɗx�����6Ptgv/�;B�v	
�҄~rv�c�����I��yxw�D<Ðv`[��Kŕ�M�{� Ɖ��Nk�	�<��#�����%�#���ڟ1�S5yQ�BB�t2�
��7P3a#Ys�W#�y×��G��3$�� �����?�Ջ��[�}0�Uʐnl�r��߅�I/�z�V%ٌ�.�S����
�ka��"�����{�:"e�*�/"���X,� 3���fve@��f��;T�����<������ ݝy���Ɏ�3te@������<t?�?ο��.�V��4�KfT�3�j��a�]��OEA_�n���4i��u����kw|ϲ�o#��yD7�T��k�|q����H	�m'j��{�sו�7x�BA��3�ޯ�����F߇��x�'�����B��WQf@��skˈ�0�튳H��[�N�F�a}�T�R����}�9䳻X���Y|Y����/�跌iy�Yۜ��Y�����I�����{���З�b�0_}d�X�Z�
�͡%ϳ6�H�'Y���p�Y�]��u�0�����S��$�\0(��"��A�pT�6�VK��r� �D�j<'�6�Ɔ-ڣ�nhR��h��9����*���P	����}��� R!p|܇:��Zo�4OԖ��l.��s���cJ�`=(����r�x����j��p������,��.��ݻ��)�
�J�R�e[af�ED��`#��|�p�P�ą�XŠ�<t�j�)+�z\u�����1go,��P�ר����*|&�.N�]�����[�b�&���L���D�+�_0����UaE�a`戻V�9(&�^��x"4�y��
���S��~#GG�.��r��)T4{1J�#��RV���h�v��0�$� ���˸���Il����ͨ�)�guh����c[t�;�#��M\_�BY�{,��ũ��D9�QuVU�8���y���@S#?�%�'~� )樚�%�C��Q���h�ߪ"k��m���=�CY�f��p8��&?�f���/Hd�m^���	C���>H��'CΎxY��O1'�7Y	^q�r����ԟ)qn��	1|��w��E�/*����q�>�U��~aV1��[�ԇ�W2e)>����Z��ڐ=�,�\#���Rի���K#,F�<�ήs��+�kg*9��ɶCv����n�p�E	���NP/Fk�U]"#���f;�W�;k��/[V��;�C3��#���J`ZJ�.v}�����fK���v�G�3�$_Pc�RgFdruT�eܟR}�&p=V�k,Y����H8������\p KZ<#�4`��!6}g9t�Ѵ՘�Ĝ.�j5�.�Sp���;�K6�SC���A\�#�!0�D�8�7�մ�(f��$���[-�s:oI�蚃��>C�����W���,\���:͎���*��̝7xi� y��8����7�'�~���AQiR &�i��9=���@��'���:��V�AW���I&�Փv��0� �6��W|a?��W�8Xa�L��E�4|��4%�Cx�yÆo%����o\yU7Z�ݛ�x���"��$M�a?v����0����K��W�8�Ŕ����=s\�9�z�ۿ�奍{㥺�~/(v��²^p{ز�QI����^3N�q)�κG*�PQ2�B�
d@��'R˳g�g
�4h���[1��]q�9���	�Y��+
B�T�m�>,s>�3K�'\c�`Zz�ZXc+����oA1���}��V~�����j�\����4���s����9k����6}9^�	�U
3	�/Vli�["x.#�L_� ��̈́
���;��|=�N�g:�-����23��.����M���"�~��B>�v���|�A"��zܧkRIj��A�.�
QFx�/^��̟D�\�䄺ԟ�fIƷ�H��m�h<��*@�ߤd��^}?ʳ�&
��������y���kQ�Pތ"�T�&-{JUc��pI�	\R�M���U�
��6�� 	p���C�8�V�;@�t�k�掆�G:_)�@����NcK�����-C�~���n��?n�I,�@��.�.�����[J�r����F�� �� �]�FqhӕQ޻b@B`��=�[�%n�5�\ܐ�Ʊ|قaeQ9���g���_��(��՜	����C�аo����S���}�n�������55���s�a�����i�mLO�$�^�&��ٜ`�Y=9/dyL��nXP�E��M7i�{�85d��Y�*;;�typ��*b�
���S�aX18J浙���38�3M���@s�M���xE}��<�i�=��Ի���v,� w���tٺ��=���#�%�^b���T��ڍb�n�4^�l�V�ߞ3�z�I��/!IIȶ��G~D/*)�9JO�·�`��5�uk���F�z
42ԓP�2����(��*=���n.�)�	.>��hπ+��v���)��d}h��V/��?8L�FO,y+�����{�����n�`�ȣ`�d�λ,������[Q1H�ʭ���FBU�n'q[ ���������1u�U���AD8�L���N�5��!FN���F�� ����t��[���������2bL����.�4���k���R�2�1X&`d�k2b��-ix�C���=�.^1U�rt,5:��/b�}�c��d��%oG��)e�2�7j��T�S�N0����Ayϧ궽0�ïAUvp,�擪ᝂ"�b6�ƍd��ډ�-U,MJ�}��� ΰsP��ݨ&�zO!��V�� �
Z��	�SF~��v�s��O��H���̿��,��o��k�Iܥ��;�J�ʑ�h�}����B�jq*^�-s��Q�r��L����ރ�H��$Jŝ1�)�P�'���p��`~"�f_*�v�"bp[|�t�.��]�Ů\��D��hՙ��g*rm��/�L%H�x��:GU'Z�c��g���%X=^�f���$�|`}~d?:19󍶚"c�͢pd�����M�l̵�s�b�\?��Q{��|�^��Y8L�;,�6�{��*�]wrVA�ף�"�7�[0�T�O�&���X�F!i�FK�R�b�#>%�[D�z�zd^Ѻ>�����p>����qyQ�]���Hr�m �4��>��� p�M�p��r���UY��c�j{D�\��H��I���{ ���x.K+aT����k�S,�hu��@��p��_H��9��"7Ӫf'����P3���Ӄ�Fu����TW��t�nC櫑5��
���`�fU��[=*}�>RK�2G���� ��2�u2���Co$g��'2�BL�>����CTD�X ̍��o���P-6JJJ��s�=L�������{lN�BJ4PQr�Z�QSEr�Sq3V�"^J�#�	�8�)��o�_-Y4'�#x��k�&jҁY1!zbq-�]ŕ�{u�h�_��ɩr7/O�L�
_5�o�ؔպ\���9�鼵AP��g�H��Y�� Nm���b����u�W]��j��W�lN�Z?�d?ci',��5iܤ瞩�?�F�r�?7<h0��^(RG_�C��Î�-�Ow2ձB��K�u?�M�p��L�ݤ�#�Haږ�<�= �4�W��GGVt���޼�F�<���Ӌ�iUb��U�D��;���(���c�"BK�]jL^�L~���׽ƾ'1?��|z\��鮂ӻ�7���`	�G�f���F^M�nEM�����Dܟ��;3�����Ð�6�Ԋ�K�3�G|��0w�G���&�ď�'C�DF ռ�����Y��baV�y�#���).���y��poKXi-��o�(������# Χ[���ݻ��R`_�T�SM�~�έ�y&�~��`�2g�f�����ўއ cP�d͈@K_�i��Jy/�J���/�!v%/�,ގ6'�ԷJpM)Z�2�]�1]��f>)1��G���ȅ�
�o؞8�8���*#C��F��wN?l Z�7J�u��I������Q�Y{z[�з7_ms�����d�yК�ݚC��rZ^�Ѹg��\04�hT�p�J ר�0K̙hm����$�7�4H�0_��3$ ��ͱ�mjO�'�j�����D��͠�&��U�!F���Z�L!,O���_t����v�Y����h��y�e�(
�K��>������;_��O��Ġ>f�z+I�� �|dNՊs��yպ��رI&H�����V
IV)Z�aeM�D�T_3�ԕo5w���j%��s�8�>B����~�
��]i�(ЛX�XD�����K�Z��{��y##R�H�K�_-���6��5�ţ��j0
-ʁ�%E�&h�7+��~��.��g��n���}5��� ����)]z��SN���Nѥ�ㄵ���d�bA_����K�`~�r�U�k`�vH&�:��9�c� .+��'��[�6)P���R#�%��+|ZI���i�Y�T*~xQ��F��=[�#��b���N��������i�[����:��De��τ9����D��[�`P������,�'������0��e{[���,[K	�8��|ޱ�=>��b������������!�y�abԹ����@�I�vҶBK~i���e��s
a�8��^QB+3?����u�b�3W� ��NL������7�$�P��V\�'h#CB'Ҁ��>�X.(�acz�^��o2d�o#���]kN���u\���3/�d,'�����G�8;me�hb��D��t�]��2tB�_"Y�R�hϹ��^�P��2bXJH��g��JkF�u�`k��1���@D\��-��5qr3ց��1�yG�*�'-lfK���n��8�keؽ�J��=+M�)����Ӹ�~љ���qwga��*ot������#�C��9������T�t3H�#�d�	���1�P��G"��v+�5E넛L"�4ʨ���܇bZ���8Z�6��W�ʂ�k�]�Z�Oی���6��@��>P�W�2�"Aۨ)���J�h�XPrp
�+�'.-]�?2�<䭞��������uϛ��^}��:��^�)5*���r=�e�1r�|�k|�@xtn.���9��u��%`>�:��;|��w�'�T��Ǚ��T��O��p�T1�ӭ�Hm"�W����}kYJT���wB3ԑ��9XπDdup��L|sJ�cZ
P����Qri��h��.S6Ba��dҢ���c�F��hG��HS��_yG���3y��&">>��3�\D��*YD$6�f��e�+�`��k9�S�y���/i�e!Zo��W|��D�*\�:�����3ԙ�����a���q6��r�,(hc�sO�t�57l��Zq_Z�q�:>��,yDuk�N��Ab:�����2^ѥhe�u=�y6����� ������!�����:���b��U���I �i�;��P�H�;�A*��C5ǟ��Q&ڋNWQ(}P�A/�\���f{�~$�2���E�[����WY "H:Z�k�r^lM��%�˅��.p
���z����;��hG���f��̊2rtϠN.C]��������_�'��e��.�۵���gUwXx�m�߈��]�\��,bI����m� 0�[��"9C-�<#��:HI�Z���9����KUdF"�1Ʊ�[���L(��a��<���]�3�F��G�38}�Ug��H��<�fU�����ܡ��6
a�`���2�"t�r�+R�2�7G� -�Jt� Fq�3w9ؖ�c�U�HJD�V�r�k�ᨒP�_v7�O+��@!�D�B�P`�a���.�(1=��O���:�XP�{�����>�P:WwF�NltS����C̶��Q��d�A�>&����ON�%�
L����M�@���3� �d����,��X94C��Y�h��Y��Bt�~{�<�����ʓҡ��ޝ��r�y�+�&@[6?��d���=��D���|�?C\���j�a�E&< ��Q�@�d�3?��{�N��������f�E�܉�K��^T�
���/y�$?}�{�"}?��Z��a6�&�OKڮ��M�&��l���n��6���R���1�6��q�[��a�y�9�q�pA���-�3UJY�~�'�f}9��d��9�V5�b�j� �`���WѿD���".���+����>~{�/%ـv�K�PP9>z�Eu��<_6��!n�?ϬCL�ֈ�`ac`O6"l4����&��,]N�>��/3��u�H+
�����E*W�<��k�|����X�%Qaczl�p�&9���$��V�e؟U��Z`�#;*N"LE�?���%�χ��
��]�+^�qB�r�0��x��������'�=��i��.�Xq�y�jЏ�#t[���9�wv�;o�0O�X����l�f��U�����PUb�ζ޻�7!L1��~�$��^�$�Z��7��5^$P���.g���nۏd���>8o+�)4�9��T�3�OU�>�r�b5���Yy�I��3%�i�'�Ҥ��Ӊ`���À�5�u0�����vA|C;I+�g�'�cn�����C���`�_��,m⮿Z	�4�~װ�(�	S\����$���Q�ڗ-���B~}�u:�ӿ��
��*Vҡ��Q��n��c��&ޭ�
��_Z��<lb��Au5j�/�w�ȹn�&ӏ;�/[�Y<������Zc�#(��h����1��ǳ7= ����V9臺��}gN�=�J6J�GT����{����9���@]�vʷ0�^i�mD��v��������v�p��|�)1<
�(�!|0�����J���n#@g#h�H$[G�����BǸ�M��W�Me!z��<���e��L�pE:�E]��xw�%~+�o�� V:%Ңs�x��;�v�}���>6L	�_2S8*��U�������+��Q�=��a6�r�7y\��m��އz�Ϲ�т�ʺ��xe�Kbn���� Yk��}Vd�zc��{���N�7g�+�:v(x��D��A2::R�w�Q6�S�8�g����3�+��,��S@�����w��G��W����I�A�6�Խ��lf�/�J���8n�]���5�<�����[�ro�D�鳒�絕�c�Kr3��~��I�����N�����".H��5D:�����!�h�	F,ۋ�w4�-��D{���uC`r���#w�/+�N�F늣�hV1�%O��}��D�������^aФ�C���y��BX�ҁxP ��mƏ�j��S[Y�����|��b��2ф�:���\��O%�N�H>R�5p����KE��R�Y	�����f��B��D�y�G�.D��~��;	V�*����zf�\��J�z���E�v���\ޞ�l�M;���胑�`�Tk�mzQ����W)y�C�+����6}0��HC������	��bV�fp�<�d�����q�������!GG��:�y�/��
J�&7o��J	�,�N}��h/a�W�]R��O���?S���\?��s�gu���Fw�������ω������R�ت}{;x��ϝ�5��M�Ŗ�*J���z�!	kԡ�8��q��֍ %G�n<���2*E��'z�����7����c���䷧�'*O��"�Ï��&�\UЁ#�$��P�����R�����|�b)�.�H�$!iۂ��ԩ�{�f��n�0@�?c���H�e�a{���2t)?;�+�Cٷ��a��+�O��7,�y�`����������h�kۆ2�WKP��C =�ERx�bU�ZU�T4��83�pL�G��KA5��҂�:9�كǏ��Á(*jZ�0�>�G���I�1���#��7���~ï%_r����,���mx����=$2A���=qe��)?dpjO�!�,<	]�>��F���1-Av�=�wD]�i�9Dm����{�g�AvB31�2"�@сy7O� ���)\J�/�����z;�q]�&9HJ��x"�Q ƢԤ�搼��cf."ۈK��M���� �Q�9�h�ܙ4;	e3�<��R�k�����0Mx�'PR6]��Om�dYA��] ��+�(o�y�b���^�D�N��ڃQϠg6�����p��ٔny*�"���Y����_�i"{���F&gi�%aюn�	�>�݈AC���.������~?�w��W�Zy� 5����2bK�쏰j	*��(�#��=ٽ(�bZ�`�9ςp���e�C�4�9�0����i��̚m}�AY��R�S⻾�GYYc��@�C���y;cאT��T���'Pl�%��]����aC�U� |��K\n_O��YON%��r�C5���zW�u�9�q�#�℁���q��i�n�1\9-=�$�ǉy�	�^��2������}��?Rau���Q_
k��ë�55�'!�Tlo�{@�,"� jP�)Q�=�0Go@2���|+���?T��Vj���&G��}ב��Qۻz��e��ٞ��?�僐p�����t���d��'HZ�#jTB2I�Z�,�~�'LˢF~Bv���<�[KȈ�M׸Z��e��Y5���neMF�Y$�}��?Sb�E��GAR��؁�k�S�[q:�J]���#�������~�zy��G�t*{q����^�a�͝���0��R�D��e�_N�y;�J������N�W�4�^�*u��{0�M�{���}��۔�ɒ�G�NL���xh^�8�lC9���*���ҦEK�cͅL�5vl�E��ߑ�>���fa�7�S�CA�|֫���ȿV�M%m�ߟ��d�����P؂i���S�d-����� e��,���ЬX��օ��b�r�I�þ	lb%�K�z3l�V��:Qcbs��gB����4���,08x˵"P\�'�6��Se]��>W胇��{��aT��8MK?p����KB�� 0���^y������q��zӿ�؜���c?h�
i�`�Z��F�@��b�_˟�X;��f�+p]���]�Ԝ$�E����b#��AOe�?���"av���uH�D84�����t+b屍�0�c��)�&�?%u��דB	���������ڑ�'�T>��v�[L[`OnXX0��M���z�@p��8�q3n����s�h,��v�	���d���n�s��~��$����uuys>��y:���y����x�oI�I@j�������up�|�[+������D�d}�Z�z&r��B��"J����ĵ�%�5(���jDAG#C�#���L��n��:�D��ު>4I�d���I���h����)�t��:K���2^ڜ)��AC�U��N��/��-A9M�b/�tq)��P>���\ $��H{e��-��9y����9XtU��>l���cK�*v����!�J��&�s�������$?�A��_�F���0��\j0:0���P~N�ԏw�&���M�Ri����m��N W���N,�E��b�2oP�:w�Q�[��SEh������G��	��"�;2�������q����`jَO����`XQߵ�R�cn7Ql'~��H�C�q���l< 65jK<�Ft�� ��0�D8��ʹÈ�����0c��y��e��h�,�,��
߳�s��Q��:1�!L<EC<�80��H�H�e�p.�_|�#M�s�A�
�c�/�,�\^���HP-��pFc���K�\!#h�)�o���oh���埱�l��[9g"�.&��!�<A���㕵V�0d��P3r���Ȧ�0G+B�
����ʞj���cD�e�~L��̱4���Ĳ',��/7�ݱ%*B��Xs��fZL�7�`���WN❿e��$<zv��7r�Ur6�����б:A�ÉC�8�>����C��l:#���y+�#}|�g���b!IR��,�(q�0�Y�Z��YC\jm��@�����x��7³�⁍���8k�#�CA?�����ȋ��+��Jˆ�;� #3���#b&R�F�����A&&:��5�����?��(�h���h��[/߹q�mk؀R�'L<V`X	h%_h[p`Y�w���}(�=4�O�P�ZZ����7�k����+t%�z��p3i�
X+z��n��s"�gȺ{�aœ�e��!dp� {��0��`��m�K ��ޥ'�*���%
p(TR���Ҝ���>�$�#�R��G�֬�H	x`d�Yd���1&����̱�����e)��,���LC �B����Dq��%��Ma�)��.�$�rf�+Wg� s[�����C@!�N�{ͽ�o���5��
&��e�#�4>94�F���%�s�v�T���9aMiWٍ��QJ֊8l��,V/:K���Q�j�lY�D񢎆��e�}��%�'�O�#����񽠾x臨�v�L5XNQ� �g6s(�����
7�d۲C0�s���{�qD����P�)�S��=�s�ｨL2=�C�l*�\��6.+��?�&9I������c���ӡ�ق�K�ĥ�_�$bςg�>����W����Ú����y[��j�	M����|';��f����NW��؋U�PA(��?�?�����_�	)jd�ЏCF��]�n�-����O�V�&�z<8�I	D@�T����p����b��i{a���#<��*�j*fsU�O�=F>��=,�?#�&��6U`�}$])1�XCv�8V��g� ))�lN���		Eɏ�tbǿW{��J�lɥP���^8�E|�l��EP��Y��A�{����LҊ�I`�@��~PDJ|5�8�k]%+-���9P��͑�wv�|q�枼�:��Ռf�+����ϖ��Y���r!���7&Uz#���*����5��A�C�!�3y�q����PE�f���U�d�`7�FL��z6�1�,R
�"��Ł�LT�_�c�Ֆ-�=*V�^��[�~/�m`2���A�Ջ���(k���-Wf�0�/�W*��(�U.'��ֳ¡dMQBcM\T4d�T�+�p�ňm/���j�W�,Ql��,��M~Ak��ۍ�B�g��.LLn�����"H��H`������}\O�Qg��*VGUњΤP´�ߥ�X� @���u�%&�8��q����W�zw���~=�'8T��0
Y8w~��������+�C����\��|p��x�g�9�H�`N0%��"6�E��hMA�Y�G4�WOyW"�9e�'���d�����a��w]��<F�ʞ�퐶�+�j�:�M�kg �O��^�����6\4_������,�vf�����=��*�Ek���1�!"7� )S���O��d����9����p	ڨf����^I��Е�]2�G�ZF"s�v�Ї�Eۛ�#f��Aҧ^.%�̞�7k�[�� Y�gA�b�������s�0�U�@�y[ �F2��Gv4S�����VP�8R����j�m�%���=�]�L˼��:�A���Aݻ8!����S�̈%6^ǌ��n� ��p9���?�i	 �Zp9x�����@/��]�D�	տ����^W�OY����ނbr������=�{A+�ٗ��0z�C̀ZC�ғW�UlTk�R�� �� H���S��Ĉ��t��,^�����9 pC�Ϙ�D���Nn�����[�MV���~r�L��g�&������p��uQn�f	�
W�񐜓l�]�G�JW�+���h	�.�
գ�+��.�+�H��$��4�Q���(��������Po�������@j9�b�k�l��X;�b=�]�*�n����^(o�ϐ���m|�7�������[��@�_��$G4/(��\O�E��"Ҩ�4�衷�N�X���>����7C�a�F�y�P������^�mn���#�	�.��8�<����S�
0�d\�v����*�X���*��׏^t�M�Z=��؍9� �Q�x�e(!�[��@D���o�+k����{������1`Ch�X�g��f@B���-�e�L�pnIH;ƣ�lAC�|n�	��l����^�;��x�M
(�<����J(�T^��j�����^	�,g��$bN&h�T��B�����Vl�}]� �n�=�
�
�38�u���;X��<_�I�^�T;�x�T���[X�]no%��a�_n����m+3�|��?����D�A1�D�����c�C5���y�H�N/��{1�,w��]QA@G�M��ۚF{5��|��*&���?������'��WݞZ�S�/��^#�ju�Q4r=q:�[a��%���H�fjs��˺x'0L#����@K� \$7��7_-5��pux�'���:�����'��y�������|���6z�$8)I��ʕm�l�8�K8����-J�4��Q���A�g9�0 @s&~�0�dþ)d�Ci�F�H?6	�
�+e�YYVI� ~���Z��05i��T�'�cZ�}�?�@각b��nM���K�Y��3a��].3u�b�cO��,���ɗ��Oqj΂�[S��r�U��Sb���ӞH����K��c~T��]�8�c�zք����6܀(0��_N��(�%V�; +n<�ҁ\P���]&yb��M�m|ݗ�N�rQO� V�~7���a:��J5qIϷ��s�f����M�|E��jZ�x{!���s�%,)	O����^�����M*VG��?��pj�W�>fi{$�Ѷ�G�G���-�ukձ��5ph�D���h�~Z;6ӌ�[�v-�E�O�Z��?yZ� )���aU��&��p���M��<�LW/���$�ٷ�߂�����=����p�-�FaE���c�S��v�f:��5����qut�&�'��1�q��s�O&&���b�,�l^Bו_��D'��X�DT�0��\S�"FxA�362��-���jrk����
U>�;=��<$�4m�]��i���x7=/�������R��R�KH[�j^V��]�!3Z�U5$0ّwݷ�-�%)�V4oˢ~�b'a�z8z���^?9�F�vD��y�׈�(Css/B�7C�`��yc���:���$3����+�i����78�:�D�Da9���ů���'�+%��Ux;;�u�����"�M*�Py��lcJ�A�އ�5�G���Fwa�?����`8�M�F�{I�"y{輴4x�G�Q�3L�#��C0K[L�b,���%�I&�؀3��1�+?x�fD��7�*�_�?��)f���j��Q���S��p��U_�9U�`��~�9Hm��+����s[��S�q����ś93��8t�Q����K����
�A�N+TT,%�6�A^3�m���'�_�d3$7r�#E6+�Mo���Z3m��t�5��E�,�M�5��4 l��1���9ݹ��!����7��}��9X�x���K:��r��V��L=�w�f9-Eb�����	5o�׃%+�| �6��f14vQ�$Z� ����q��=�<:�24��T����x�{?��������-@�8�Q%p!�6yʦL�����ˢ�pf.�夯+��Ql!=��O�#E��Ϳ��U'4R~���U^�~�m1M��$U�'n&᭷�K~��h#�0-�����W9Ѭ���r�TʤS�b�h�ˍMb���d]����=a�,ߩ����>����A�,'��E��$�."�^3�j~�I��~l����ǹ���s��jH;�t|�8�g�9�R��'vEU��2U=�}"�m�o�����<6�3y��}�Nh�`L+�`$����8�pΒW3hE_��Z-y8�T���U��W�^�n�'�45����̿W��S�:���ph>7��Q��潉
�Pޟ�$������������1�D+)Ҷ�;�nMh�(m�p�[~B��ר�m��^δѸ��i��s2��J{��r����h���X#B��J�o/��;�ȅ푔,���=b����}X�s�k#��j����M�1]��Lc�l��uD�.By���v[.��� &��>��Z��F������E#�M�z��r�&��� #�j>E�?U����ݪޮ��9�.��ɕ��O��Ń���1A�@���p� �eO���$��_�y%�,��*�>.�M�	>�����Q�>�� �{�!�!H>v��^$���q֖���R�Ð��(߽#�	[*��m���Y��d�C��ȼs�pfu|<L0i1䝴R6�����WIø�g�R`GR7݀���j�������r��9m��j�=�V��YTж#fo��vJh��M*kٯ�&�.H�zm{+��I��2Z!6��{���L����RTT��_tW�,g��1La���)ߝ
��X�kQ�]���%sEV�y��0sP�< �*���պ0t*��U�T<r;XGІ��^�[�����$}>F��V6�o#��O�īA�����4+\�GM5e����ފ�ZS�,	L̊UTL�QSS�� b?�T�[P�>�㦰����z;�����
\>�֪�C1������z@}ѽ�$����=�h1����jtTT�@��& s�I�@��7au�,�*P��p��ARM��^�7}|@��-=>��	^�\�c������E1�x;����²>���Or���U�� yMV�`�)5)�!�����P�;��X�A����C;:����Ji�S��rW�}9ܫ\��%h�%������J�e�]So9�f��\F�3�B��p��#N��e��f�)��S*���b�3�Aʍ�B�6W�F�_&���i�4Ѹh_'���ew�{:��;ݾM��!u�;��� P2e��%��8(.1*����R�E�g�Z���a�ҐU��{r�-�F���$��L��g�V���gLIx���w��7|@7����n���I���-mī b�>T3���Z$�($����L�_��V�Y�R��@i�����@�=�
E¶��e*��;}ԸV���g�؇��*��O��"0۠���<ED�##�ү֫�6��N��n3;�Mk0�*����H�H��!��mԢ��EItG�>��g���v��8����u��k���3���l��	�ws�j}��W����XP�I�TDNܠ�r�J�Q_��MH�:�$A�C������;����CF(*�����z�y�5��d�;J0�R��yxF�����ZN>ɤ�����T�dH���a�%���V����.���kZ�}��J�5�?dm�/�,̂���6�9��{�@ ���lUӚ�=�䓔a�Z�zo%���	����s�s=� ���:��j�`N���H�	%�*��(���ȗ��$��+b7�4�A�HV�xt�U�ғ&�d��o<��W�'W�#��ң�U��4	��Z�������{���Mo�I��i �b ������s0�n��{�&�YvO���x�
W�3��s���G/����l�d4-[]��t��&ΣT(�)>-�z�cF�;4'�(7���o�mJغ#���<	�!,"�2��)�G;�=����$�6�*}���O8hQ����0�^b�@n�����zh�w���j�w�)Yd�������w���@l�%Ա���n7���f��j��!E2��μT�Pz����8��|�5�_(]f����:�F�\6�c"қb��^JRZ#,<��̇�;�P�v?��]m�t�Ơ�%�oS�0�w��)���$[� ��T`(bE��((�-j=//U�uH��@h	�}ݳg��PP�9K%�����wO⎯�q/I��x�n~�#�W�|�=*���B��*��Or��
5�D�G�c�����z�]�s)�狊'[o^l������ܻ�����E��� �5��~=G�*��S/�x�T�����Wz���Q���ՓB��&\���Ve#�@��QWS����_/>��]��9@���}+r�̔���X��-�>F��?��ҋ�Ɠ�k��R���v\u�W��~z��ByF��nBt�ã(��E�5�,�����kZbZ��D5�~l��^�("�>P�鸚;�qy���Q��#A���9����(rt��g�~eX�he�bw(�㪮�\'�%�;,���-����b5X��Ҍ��q>���>N��~Dt����C�[�uD�%��`۽�F,�/�W:9w��;d}��A_m*N��m�|�hߙ�N)J�	H���~G��FC*Ӄ��]ܫci����J�h/�[e}CQ����[3C�R��Ԝ�W|K0���b�!���������}���V�@��"�
1��~60��lj�A4�>rH}�ZN���&�-�-#���ՃZf��-Ɓ�d������.g�g�(�/R�1`��L4���*QZ��a[�'���k����Fb<l���u���:XP
G�J��v�0@�=�Z�v��A;���w��ɻ[��x�4�i���h���� �S�,F��.�}��e���Z/����w(��]�#���_ۂ�1)��E��k��Ux��z�@RR)�n����u�%��j˫B�U�JO��&m�Qh���}{�=��
EhF:����.臔|�i/���ħJ��5/�0����W6��?^-�!T�avhg4��0bpq��7 ��|
�j����h��Q�l�����:?"3)��$��{��@ɣO�����g@�h�qp�Vi'8�!D��4������9�7�/��I����u䅽���2�f�MN�coGV<��p�t�p��$�y���WΥ>�e�M�Nֳ�� ���}�Lf�̇��̖������	�[�*%���%��n��
���b�*��1ò����	��D�6J�z��q'�|,٧RF�&D`[��0��\���W�U�)�?[˼�����e>Z��=5H"�(D��|�-+aU�NΟ��r�ƈ� >����K{r�pD�r4�̫:��ڝO���L:��w���v�Ρ���hC�mh*C���s/�we0�������r��CAci��NT����}t0�����7Z���S���x̌�B=�E�d^��_T$i�1�bU�Gr�:)�>��7	�@;�!)Ŵ��W*iC��X���wu`�
�Ib�%L0�Hl�[HcOBD��g���VJ5�a�J����F����<+��Kt�d���B��1���M�D����6D}��5��+kn���Ob���J'�q-k
`9��P�����e�w M��������IOSF�D0A�
�@A�q�/*A}���;m��)~���Pp��1���S��k�#BŌ=ub#吂Ϋ�@��ݸ�f����%��vby�z?�M��NE����(�m������e�����7}��l���|���b�����nn?[��o��r�B�2���\�IZz�_�H%�E� �� ƈ��g��H������������-o��JɄ�.�e��W��%d6B'�I��ZQ��{_1z��`צ�.Q:��oF9���
�czv��)m�:�$�����f�cyb���_󲰈�A��bk���$�f��t�Rjl	�v|X���J������a���n�{�ziF�ͦ����-b��C0�l�X w�����m��d���Ț�!
.(0p�eoH��Wy����|��PA��&�hQ~��������n�a4G��;0Lbm)]��v6�N{Xt_Gi�;]Ԏ:���oG���k�;?���D$��.A��J��h�=n�Z+��<�'��ea��\��� �v X?���^����!쐫���^x�vx��q
z�RV��+o(��1,�w�I�:�[����r��[e�'���D�:W���Yܩ��Y����[�~�@����],�|H�O�%��
�v#D�8\u��<�@����&h��p9p鰯�:��+����WCs(�����'߻�JՉ� p�e�k�┢�i����% 2y��m����o�H�(:�j�����LAhNR2�叫�Ot�+S��D<j���j�w�l�i{QP!+����N�����i��/�=g�&Q�>�~X�8�ov]9֗�đ�-����A,��Y�˖�o�I��h^R�~V;	��,��/p�&�aQ�i��`���2[w����#Y���Lxͣ�J�s����D_Y�� ���J?��N5�-ŃWg?��^��@0���kvxuȱ�o[%l�Ls��)�a����9�Yiҏ����_��@�"à?���ŧ��T߫�?-�l;�3�)�W��Q1�(_��ŋZ��E�(;�牵d���p������W�=	�O��2�[r����d��h*��3yIg� �=w�����v/�( i��N
�J������wy�p�5"/f5��ٝ5"7������Z���p
4�������U`�$ ��)6�����a3�ϡȴ.+�����`������wjx~>��}��HR���,�܆Qb�u�	���w������.D3Sc�Y��!���U#����^k�dXK��#�6�	YR~ >}P�1p��ln�\���***/4�>�����l@ �#V|l�~����]aa��3O׎V��u�l���?�w�"��y�b0l�_���,�ηR����\���hB_�>�E�ʨ@�\1�d|��Wf���G�c�<�t�z	kuQ���.ʋ�N�C�|�Iu���\�qڧ�0�Q�k�4�F�$�!b���y�WЙ��Fj��O*e���I��&��#mk�e�L0ka��'�[���WPhMO<��X�I�[c�j,��iD����U*xo�7ɳ�~G�W����/+ao�,���n;s@̘�i�V~]��k����F��0^N�Z��`���-$~� C>0]�7P�4.�(��M��=�3`!J�=�v�F�k,�tMAD#�4��������y5�RB��,�WX��]�a ���T�C�C@������R���qT��h ��"Ā(�M��!)3���1�^���C،�r5�4��w�21H�A��L��W9b�m���1(�`b��Zl��3҇,��cGm+�(�
��Y��.P���i�s�|u,�P��,+=8�o�oKy#�P*^�	�w]�Ѷwgχ��Y�k��"јi�~jc��s]�{)H�3���eC@��C�qe�U�^f�G��L1�?~�?wobj͋w�eI?c�fߚ����J]�6�K�/������UZ���]�tn��jW�����y��P'���r��V���Ɛ(���F�����R��b}����G4�3�8����jϸq*$w�0�?xI�|*i:?^�ca!+qah��(�A�#L��=�����-��Z�t�/�/���B���v����	�Ǡ�5��Om�䰄��w>8Q�[����\$5��s�'�����BBq�+5�%�GLkQ���:��91͢��bQ3x���RO�x�/��5`^HNw#�Ϸ�f�4ƄfE�e�\�.n1���ȥ�X�*k�E������w"�=����� ]̀�J��K鸄H�CVm���'�����T@�� �,��G�w(�R�t������2e��ɘ���2��!;wbs��Dn,yXŰ���=��Y݋w㝆_�I'����b�'(�dB��ZV�<�US�o�cI>�o���d7��Q�&�B���-e4ƣ ��n���A���%ߍ�4��#���'��TM/�+��Ν+aX8�E��q�� AmL2�=�^� �*%'�q��m	����� �f���mh��h��3=ٗu�}jç����.�P�K{���_�[��QC��Mz�;~�f������b���r�˵9t'�G���LT�+��\;t䱹�^����i���#�<<Vo��|6�^���[U� ���R�0�!�n�bIe�c�扬^3�~6){��Ņ�u;>�C��>�i�߄�@�1��jՉ�t���H�����f݄��C4c��d�&Wߠ)�%]���1 uckP?,T�����o�mq���w0��-	K���,��Q����i�\<��P�i�GD��-~.0���h����ī�<�AF����g�8�~~h��;�Y˨��ay7����Qc�7�G�(�ս�=J>���#�t��P�@��-��c�T��Z�4��$�cQ�^q�0�ʣ��ё6W����]'�^G�����������TP�a4Xe)L�^%p�I����g���9�U]8X2��8|��\���<��]�����"�c9�d�r�61�KL�w����X��d�xu��G���]t؎����X3�y9f��K �B?��/%$��Lk��x�q8[n�~Է]*ˁ̘��`�z�d�>vA���,v�rJ�H����d��fl�DÂ��]A� u��;�J��H�R����z�3!fů�H�#�n�/A���9��E��-4j[�h���C�u�����
����E4@��q+T��
�+�
������~�{3)��]˯^�v9��3H������o��"?�S~��q2{��A5j:�� �z��ٳE�$�<f时�p� �H׌�YpKB�rq��roY
���k:	��eR'+����|y f
�T�*̾�?���Qe1�*���91#�������R�RG��o�`����_Ⱥ#�w�BY�X���6�6�CǇ�?��Qv���z��h�ξ�80���?+|m}� >W�é�@�bb��FOጶ+G�KD$���_��j����߃�˭�6�vH�ķ��V6+�{#,�;�T��m��1S�w:X������6��$u춐��e�uW��CO��3ޮ=�0�{�9\S��^HQh}�f�����~^ŷ)ށ,�vev�+��v���!E��*�|���l�¸��S���۝W�َ���x=�U��ny�껛�[h���/���ź��F�_�œ>�"e�r��2$��Q�Ⱥ�s�����r{X���'��ub�c5VԱ���"%'f@�ܖ<ܤ����`�i��55�/Y��B4A�f�E�퐠E�&HC;�T�@�d8X����|�F���i��� y��yf/����"I��Vy��rZ� �]b�h;۔"�jx��џP�I)�6��͘T'��T�x�dzѓa���ξ����|�ȹ���U�{�l��ΖV�'k�Y����I^��U��-{Œ���`ʀ�`2Q`Bt\��0#�`�`#���2,�p�y5��]�h���&�"x����]�r�8�z�0�}HRF�����[�&1��K�	��R�(|!�Y������bd�L����)�S)	���0����_���ךt��@fd��&+��΍��g�L=Q��xR�[e��-�W �2�[zD�d��B�d����s��&��&�D�`t�/�����6�z���Xw�kͻan
��<���~?�QI�� ��K�*tK�[��$c�@W~��2y�׏��ϕ�<���&��"[o�Bѕ�H�~s�IJCe^$�B�	�w���=����q�|s���a"���y?�g�D�:X���6�yT��㳨�،�S F�x�YvqXLCB*�_�8���+�5v��5�r"�Gqǜ���?�J%�0�S��@@�L�S/HB��s�n*��h��t�#�j/���hk?�������N��w;���:�m��ki����;����^��Uf�`�#�]U��-�N��!?�e ��#mLN��/���=Z����|xæ7w	���#����3&��d"�=`��&N�_{� �s��h��:?�0zS�9��u��5�{i�N3������zb�1�D��'��[OE���܃���"��}��U�i��4Da@���qTd�a��g(�%�H��?ZX��=��p�t�Mv~`�h�B�X��Ff)�M(�qb�m��V���s�6[��ܒ�Or�Gcq�p[霵tn����Q�Q?��E�=�.���W��uv
q*B��&Ǎ�O?Db��Ѡk�r�H��+8uB���[��T�
�W�`�W%�SÍQ!��NI�|�/sF�|��co���]���Gv�7��]�F�ʙO�<��Vu�+�=���>5<  9�yp">+�h;�d���#��������"o)��|(�$]k�$��fQ7i
^J)-���Y�!���nE+X�ۃ�E�|Ҟ7"�|�pS�����[�n��=����$��xVexB�N�n��;oЭ��pH�e����7M��|�{~��{mh�}�Q.��4:K������{�'�M�.���e�(�Qxo����U6^�`wz�CXYe
nC�%�nk�׈e�P!���1!��5�Y�	�y�MZ+O�i|���v��cZ�Ł ��Z���'�"�qm��.R�����1�7\i�hU:p�d�Ғ�1j�Z�z|�41�X l�ɥ��֗j> ���s�	�[j��j�H�B
3��oݨ���f3�ԋ���	��ӝ6��_�s/f )���g&��V�q_.@@4�K�k�.��lM�O,��G!�DVoYz�5����Y�Ok>r|�eA���c^�<����6?X��8��0S����� \��x��Xzt�>�~j]�az�d�Ɍм����7!�~��D,'�� ��~���<��c&-l��i$G��H���:�r�Mu��(�k�Xo�c�t��J[�9ռ�Ïm*���R?�{z1	Y�8�V���(W�y��Ǥe����_�EM�*𕧫l�:6u,cX�.�)"�jI��C\���0�����r`a�!cަ�>~��/����6��a�����0�{�J݃���Q� �xۯh��z�	w�����5,Ő�i�0�2��;�<z}����֡j�R3�~�Ĩ�D.O���ަE k@=9�C�v��M9j�����]n�	�r�0�=|Q�=mԱZg� �Z�R˫3þtV�Z��ٖ��9���� |kw��k��V=Ӎ��G�^53��l:���.K�����i���;��FE����p7ɟ�����J��)�P���_�ɋз�ə���v��bb1�Y)8��!GC��mr�;�b+���M��j���c��
�_O�c9��Ǆ�G��#�"�fE����	IM�������� 9�Z��lӪ^�������x������w����'<����!��ʹ�W˟�.�`
dYX��U�S{���X�2>E>�Vo8TX��\r��8��s%��:��j����	
��m�Q�^������ +)�g�&��LIe���V�ZQ����X�Va��z I���K�Zʗ�����SNb�&N�fK�ځ�-d���|m�Vs�O_?}�1��Cijz�7��
����%��B>�Bp$���#P�[$���=҈Qi�,`ۜ��휋�Y�C�2�[��&�~�u�y_\/R	�^�1"A�m���#>�^p\1�R1�D�M2���v��4�>��,�� �u=%qh���=����L�
/��tQ�xy��DO��CSq!��H�*��a�������t?3X�	]×RL���AC,��D̖�9����;�,�����$֣O\��̙A-�xp���d9}3:���Lgƻ6�n�@��#��V��X��d{ʝ;�rbMD�Zg����pX�.�V�{����Yv����κ�sƪ7&�*�N�am՘h��-�Ka[C�-������4�_����%Ǯ1�nIp�}]O3}�#�'�٠j��I��e�4LT���	
���\�+JL{� +3��x�i%�Z�|҄�C:�E(��xSU��)�!;Je�m@'�6�N����u{��˷��)�(<K�4��T�����DM/��J�C��f.T(`�w�ş� GU��aN�x�-H7�Me=֨E�C7;���J�;��Q�i<ˈr*|(Y��φ���җ�����ka����Q̙;9wƧ�Nȥ�3`��8p���j%�u�OX]�$��?�A*v/���_n^�\g.�@1�_-�9��w�^:�(�/�սdeU�I�$�
���Of[��MH��/���CN�n��Ǻ9w^o*u3���jS��v�г�[?jv\79�W�F��Ώ^��Ʒ�L�t���P��!���3p�=��}�u��5SB���ؓ�\-37.��'��ߞ�)9@F�}dȷ�*�54�g�ێ3[C�.�����(C�8��|�� ��������J����t$�K�KD9��Q��>��bZ��k>��l�}��YdsE<{U�q!7�tFUc�B ���=ؔg�S��@$�ƹMá�Ƥ0����P$�Ż�s{G��x	�O��{n>�2lzČ��xq�u0)EO��;�P��٫4�9��#�_0\l_2E_�j�;=�L��x���m� *��7.`.����~��~�	���oB�R�/�a5���gh��XO�W̡T�?�|w[L}�2��	;R\���t|{\����JA��ȴ��1�����wD:@F6I�Q8���c�.a��w�O/�*h�?��S���A*\�L3F����أ�� ϵ	l�b1B9���q�?��b��Ͷ6�]k���� ?�D���g#)���_8U�d~ۊ4�Y��[�!��_CZX �!�(��#>ǯ,�ҍ�,�_v:o��v&�33m�'��@�������x��wŹ 
�7z�\�ʻd�#�#���YͿ�k��4�RrŔ�?��ul95�N�fT��+ \�W�Nd@��ٚ��P�'�&-�TE��%t�a���$.������2�6�컊[!��?�h���׏���9�� Ő����R_kz��Ε:EV(׌�Yq�Lx`OA��Oy��������WKYjX�o��e�#�2��� N�"��D���IǺ#y�_�G�`��l&(՜�m;��coW��~�L�r�	C��X��/�ː��vѫ�g���n�D����*-�y3��f֧��6F�cMBt���;�
y���E���*�	gS������[j� Î�۸y_dʡ��t�{k�!��������tJD`�X�_���T�EX�R������x��rx�*���}�3�z������gK;��8�+F�I�ql6�uFui"�<ɕ��,�R�{���A*(���0_�LV�j�ߧ�Zۻ�VI�n�{��d$�j���o, m!^~q7 "��*�9�2�e<�x�,�y|쯱�!�ly� ��8�L 0�ѫ��<�V��RL����=E{�����C�`�x4��c�33�j���G s�.��Va�n�awp��#�L���/ƦP�N�Y!e��#�����T8�^��������X�#�|���v4yݕ���	��?�ʿ�D������fʃ�y��:�e�)6��Pj�1�+���z��i׭o�Ox^�žk� ���%$w��:��SB4a�d,w�?#{�ϬZؕ��A7���� �uӴ����wN�4L3�����>���f������JT����jq]Wۺ��m�l�&-����?�`GeS�k��>��g�r�(�8lQ��/�D����7�{y��_f}�G+�b*�Xx�_d�>e��� \w_U��A���" =�.�����B���:�Ȩ�Yjs��j�+�7CR`�2l/�ˢ�G�Æpp���м�>���?�5�>!��?��Z��?4�? ��S�ܷ���l:�Ns����B��<�S{�g1�ߩt���-��7����������s��v�W�}�}�Dvs2n, �����r>�;�7k�S������=��PҴ��0!���$��fBZ߫����(*�v�J��a�����O´[h~����rll®�~?RƦ����L:�O��Ud#�~`�Ւbұ�.�T�/�H4��Fos�l}���ð�P�z,�(��#g#�H M�Vi��b<�e���7{-����H#�,Y�j�<0 ��|���a*[�ݰ����:�37T��Q/�����Ƣ���g��Ou�8"8e�1l�tJx���Z&�D�}%�e.�[m�֎(��a��ښk�>}F�
��d���0O��C���N߄j�|��ߦ�� �W���W'c���ے���y�t5.�8���[+�F����Կ�A���@T�@�;.!P�"C�ʿkFa�H��"Б�|�-}���%3<�,��P��������_]^׾
�I�O��@��,:�\���H�8�h������D��Ő���V����L�hHc���(䀜7������O�7�x[�<��Bg3�\X�a2�.9yU�~�3S�{���p^�砳�(�#2p#ݖ�p(�]ċ��#�0��r�U@��F�\ͷd_��X�?�L����5ҭ�Y��ժ�0��֨��/�s�?���A��떲}w+"�q���6�I�����<�y�����5)`𺱙y$���)��B�W��=Ӥ�6�����Z��r���K�b�"?i?`G�0�;��k�_C�`X��[��6�.ϊ�X��� ���	�"w��dW�>�����-3%D����03�W.�0�D��#uд0�Ś��	��,C�4�_d(������l{�r7sQ^Ș�6`�� lm����W�'z�(�_+[7���ir�*0�[E�ˏ5��_��ی�����߲Z)2�vaw�%���=���::��l�ob��g�.��f��jb���k�J��ƪ�\Ş�/���d�<w@r��7��&���=�T4��`H����3��k#4��
��ǈ�?����o��=�����MB]w�������p��V�я4,���O����&8f�oj��BR�n~I[[��'�\����2��9_�@�5`.�W8A�ǫ��l�2$Gg���2֖�J����kkw9�W5IP3���%�?��A���e��� M� ��X$��4)[r���(M ���-�,Ǯ+ٷ��Ӯ~]����?[J���[��q����'3~x�Y��v���Ǧ3P`����<��LB:�ezd�y{����o�@>��^�*��~�s��J��3�o?��'���]�|��%ʇҘ�>��(C b�r>��ɲA�k����L����{Y���X���rm��Դ�R����%ZT���a��B���k�i����<��<��P%:�Z�{^����N����S�ݽ�=�)�{�ˎۿ��;�x�a�i��<Ѱ�|1"
^�0�|q�}P0��$��M�381���\�:p������P��?[5��9YX��O7ƙ���b���Y����W�
qw"č�Ԁ�+
�a��Y�e~����|�̈́��PD�����k���t9�*�����8�����T?Q��^��Wzw������3a��P�����K��� �ޜ4�q�:�V���PES\}!�5,���"�5j�
N¡e��ŧ��.�s�m��.�/S��'b�}o��t0�@0��SVPP����"���	�O,(N�@�2uo�I�2�B3q���)���7��D���^�NW��`K6�S�/�J0W�_(/ٍt��n��`(&q y�U�I�L��o�V�eZ �&��K�z�dm���\��i�q ��/�}����B�_$�4�(*��A����h���>u����2����&S���L���FmFc.�b7a�םĸOR!0sMv�4?��������J��������@��Cu�	���$��+�,�Ѽ�l(��,t�nsK��t������NE���B��{!��i"�k�F�^>�8Uyc�ip��1�8���^F��A�b�^��W.pG�n�1��4�mF% �Ӝ�K�M�YR��$g+���F����<�NS����ri��{��K���I{�8x�ৃ���?��I/-���^���!�Z�����m���@$0���F��4����U�!'ɬ�:��TՐ�z��
����O����A�	^�ߵ��XD�)G�G���g���~픑�⮗�.�ڊ����6"�c�vC���ѷ(Q9��r�D\�R�C1I��� ̛��BuQ��P��E�RM=r�օ⠾ ���?֠��9qA�h�(N,"3��'[/F�7*�GD��Cn�����N9�\�53���aW����ԓ�Rh#�E��������������h�|�\y{q�~�!�(1�g��.���(�AC���t�Z z��1�lG��`�6��ՠ�,V��GY����;��Z��@���5��ǔY/$�Fϼ?�R���F����n�=�Y)��dq��%�N�0/H	�SȯdAJ�WO������SEnR��g��*ͽ�s��Ύ���[�ߵx���M@I5�s�����7�@I��"�]R��ɓ� �8��=�=�Gu�;�E2�<k� ˿$0;�4�����\�/m"�N�;r�N{�,�:BxܔK��~�~s�0�0x9���h�2���^oΑy��+�o�����g'����=LM�u�f����U��0�~51�}���0$Ys���QMg�1�1�0�s��B�����>-�]���B^n��C�Q��a�u���>\3�`�:�uw	�y�K*d�ʊ�����TH�+�ۃ0:�ޥ�]m�+A$.n�*h]�+�3�d�g��J31��u�=�����*���]� �',;�^A<Tc�j5H�F��em����T^�Ñ�"^8�Or���f��6@�j��Y|m�=<L�?ء������u�T�B��	��t��Wu-��ԥ 0�l�;��4�<�NT��߀��;X���������Hoo������dog���SCpC(f=>�O���K�;������-k^�W����d�Ռa��9�#�6�q���2NH��t�{���'�FNiE���f�f� r�&ޠ�X.r
�<9q+l���?��:�r�co��?�S��]�^4�+3\�NAՌ�Ѱ\�o)�@�#�d��D�m	j�y��O�=v�<�2���;I�P��/�u`�i��Qh����c3�tUy};̻��m�-X���#��J�Zu`�8j�:*Ȁ���o������u�d��lX�����M�ֻm��tJdK����
U�Ii�EfT-0�uRg�wC%.���.�G;�Ŧa����6
��V�f�͊wGj��*6�E0���o�JZ����ɝ#�3S97~*q��bi&C� (� �H/WN�y�L]SDo�����yvo])�J�HEȶ��(�p�}��d��r�.o�<҆�;��$����T���՘������jPC0��6��FJi{�[)�n�c+<G�P���p�����t��nX�eY=7w!����GJ��=n��TZ'K��T�X(��ml�H�|gd���g�7�z�|��ylK]�ء�Ȓ,	5h���/ŬI�7�|<X+
%�hc,dI���.
���6����$�NDp؋-�����tn�W�Me�s=��&�[��\a��3I�ƍ�g�����'*5H?��ap�V�ͭEy�0�Mp�VZ6�es>ɧ�]�{��fnE:��3��&��H<�w�.Ҩ�j���Ef68le�;a:�I��f�M|��L��,�<�q�b�_��8�7؇��6��}Rn����%\�z1�`�Pq#�[��q^�[%*��(T�����k<�຺!U�c��{�Lj)rm��<�3�M|-����X���s�"Q�\�{�!)1���;�G�4���1ڄ��G>s �pj|_PG�KR��B���Jܛ(�lM�/��#�m�]��S�L+t�'�O{����D ������Ɖ���zDD�t��������r^������o7H*�5�򮢃QTR�ߤ���q��X��<���`�%Lu��JFdc�
������o�rQ<���.v�d�~d6����d��\��R�6��,�h�G���c@a��*�bs�ZVI�3e�CMU��ʟ&j��O��н,��=��]݇c��f�3F�uԁ�DY�j�JD���&�a��G�����۟�P�G ��Z-����bk{g�C߷�ے)sb�ל���2ڬ%�{��]Z4VR������#+�`8���N��|��28\�=�I	<�ŌC�����!�e��J�@�C`0���e���d�Oy��\�]޷�*��M�Y1�+�tZ��=�^�i�U����qx�Y��[#:�3Ey��K�Ua��#������]�X@-(6��7���n2���y�3���kyi�L�^�ڋ�mQM��s��	�s\(��&ǂb�A��H�����-�d�ֈ_x�a�Z�B�$�^��W��($�v�7s�q�$+|�W�+�3�8�}7����#ގ��Qj_��h����h	���.�{Ͼ��1��,ˡ���W�� �%�b�K�l�M{�K�>���_g7�XOe���|��`�v���zr�[���L�[~�a�S�54QM��.�E�:�����s��\� i��2�]��P,�nR��ތ��1�լn��mFT�ث<��Y��=.�1ٔsX0�-�*�˭����p���λ�g��2���m����|��vr��B*>+�w$;�X%^���q��i��<ǩ�utD�XƻA������6|h.[Fk����~,�Q�NX=�۩ra�ϳ�(���xt@�pOK8�O8ң/��纸�_�W�h���е�T�i ��w:V�l�ơ@����#�E��+�B�h�#l
��ht����8qcNiN����>���c�n@��bz�0���aEM��Y/��&�M�5��Yob4�m5}��Ր��R�2Y�w��6`�M�����q�C��\�h#�զv�@�M��~�%�W�������N2&:L%�0�tO����n�m���v���l^��M�\&��#ZAͥH�r�W(�T�u�'v�����J���Ҋ�����*��(\�V�uo�!b���$���,&���Q�砾���(�l�h+���χi3_|��ruy�����z7d�af'�᳣�'qO��"Ҹ��a��|˶�EgPW�ܬ���!b�����<n�"��xr���H��*���g�_�	p�K�I7�<��!m�o$SbP�S�����"�u��:�H=ԍ��q�w��<ȼ䤟/s�+<�PGxϞ]�9L1�:}s����-��?����8F�d��i�q !�6� �Qn���� ɡ��kD��I&s�4�|�B�Ф�� y�3}�	;]��@�
G�aH��Eb@�"���]bE�H8�8�W�i��Ǌ�9�]�{w�45��d��^,���uN�5x!����5="K���g�t���u8-�`5
�?y���~�-�;ޭHa#	�1���/�&E@�f��
�B�M�7��E6Hd{��(f�_�� �1Zݰ����I�T���A�М��r'����#�4��v(�h�>�R45W�cl~�W}^�����6��d#�7�d/uQ-m����n��t��F��(�V��D�������`b��ճɴ�@��M#�nF���cN��^��XpV��v��j��W��/�|]w���m��<h��*1��X�g]�*ϖ��7��ӏ�[��2hGM�%�>�S=P^p<t��e�T|�Zp�/Q�Ԑ�+��kA7
��"�q�ᕝy-b�PS��Vi��Ja����Ji+G�����ubӜ6��P�<#��������/?���J�V��>Fv5���.��nf�����6���6ϫdI���`bH-�ߝ&�AQA�:xW�����Y%��_��i+l�hbCE������ ��9#����ߑ3VZ�b4|/Hl<u�T��'Ϛ��ԇN͎cc3H�0�^$� ��<�	!���V_��ǭ��N�xKb��/tJ��*@[�L�/�(fx���Eq�Q���R�f�S�DD�]�������r`Up 9��#�5��h��>*��oo�	����c�)2�N/zl?N�i4C8���@����_N���z��hTV���E2����k�?ÆS����X�F�k�w��t���,��Z��`EM=�ER w�"۬�`��x�jrTc<�z���X�������ϗ
-������a&��e�	0��a�\-oa/�����s��9����C���-3jx�
�6,�6���й�AFn��=�)a���c��.G�x�R�H_.8�p*��#q��QT5���c�>�0�^^���k%ԃ:'h��`��3���Zj�>۲������:|	X�h
=���*�dPLTI���d~s�
�:PV�����ۧ g9w��wA�B R ��G#�o��l�r`��@�L�e@E�������o�I</��� #f����Jlz�N�âר�ỻ�2�T����<"�6�kF����Z���w��Q���׼�%����H��ϸ̾� ��)�H$�ې'ہ�7q�룫�T��q��/@ń#E}V3��/����T�}Y��-p^�L��Uh��M��Z��y��ӯSbڝg���Q/�Mg��J��-�.|��aa�=׵L����G	��b�>���x1R�W�k�g�)��"�qiw��P�n�}rut?{*�Y{���_X��j��M�.�1�wƛ�s��b̥[a�!ӉX�u���65�;&-?Pl�L��M��vwt_<�`?�b@�]s9%?�NmĞ��	i�ʹ�ل%1 �9����I���hj`��/|���.���`\	!6Jf�*D��3%9i��"�!��?LbL��`�,���U��<�mV�K��l��viR4pBH�~��C���tϋֱ�t4��i�'^f�>�oz�B���^<�K�z�xI�����N���sD��DN=s囕�%�o ��Țp��%'�Q(�o3+��WH�m����Χ���G����I �Q�{�ಘ�x�kZ5:V'��ol]PL��i�J�o���Bx4}�Ȅ��<���K)�
=����8�f���n�ݗ��0�RQү�'�!^�j��ڼl��D��5.�� �K:�^~W<�od��"�����I\ �Bju���PV���̜%�M��_+:��!�罱]��� �T��,���υϪ�{��W'��y�&D0(������^�&��<�`�g$f�XOS���|��V �1>P �~�R!����97��o����~�Y�{���5p鐹���ÔV�7��]RAjx�0 �����/��j���C-�$y;w�!����b�I,�QY��h#k��O�}��9��wD$�W�v��`��d%/})/�=|�wb���� P���S�0T�z�P]?�(���lԤ�� 7ZH(�O�oNqr~�Ӛ5F�y�ƛ �6����޶��e��W4@t�	��a+ n�������e�;0!C9��B�8ݴF~�����7׀#�l�ֿ�#e�͍���JIg` ��&����T�t=:(�VGrC�2�Q�d8��d>���)@���[��G���hX3�r�N֟�U�$ptS���CX�@���ż�����J+i�p�SP�6�/X8���o�!�5(v@*���==���0�`vW3׮����h�����n�k�f��3�\^eW��|�hnUzЫ��/��]��	�G�{-�eE7��Έoda�K���`�!L���{ɧ
��ȅ�B����%�N�딓�A,�3�]�A�����:p_/*)���iIK��H�4�Gm����۔�`I�Т�N}�ݐ�;�y�Ku:|4�x��\Qr�l������D���Gf���`�0���(�e���+�{|w��H�j1�[�m��٣Df��t?'�����{��qg������_-���sw5a[\0�l%��ލ��?$�=9��@P>����O3�if�f[֨�&\�͙��B���L�{K/!��cR0�Ơ�j��ܿ�����7�}���TMaM^�0�_���	����)�R�2�-�o[e ��F�� ��g��Uz@�C�%�R�O�}Kv��{L�!�+�Ɩ{5��k��h��\����9��Aϴ�uh^�/�-��l�,��X��!�#��+��������	���&x\!�Mu���7��!f��h)�m��)�}鮗1=�,�k���8]$�Lm��ϛˣv��et���R�J$|\�Z(�o���ɣ-���`V=�s/eۤ6���?���ߨ��$��1
���aK<7�9m��
��F�����X�_ �"��4��@U���y�f=��xAf8[�p��D�XYp�%e`^#��Í����n���}�\l�� �wB1���^:}x���&p��Φ���<�)D]��J��t�y8��7mZ��QW��Q5��ӫ��'�z(:]���bݣ�u���w��%�eh���e�����l�E��ڌ�ǧ�ڃ�r�(��u���K�������-��d���w��F�	![v��K���c�":N�{a���߬��T����3,o��R���~%����3F� �.%�0�;�}�M�!�����^:���X�
����Vm��Q�n�c#=�u>�˄%��m�j�V�[-��2����1!�d	��Y��5��3P����ši:j�Xq���.=���!���"f�!�fŵ4�>:���F�(F���-���"YIj��"���݈Up-Ő�"����Y,�r��|�i�ܮ��˧��۞��a�9?��ؙ(NEI��G���s��G��<�]ĩ���5�4���ȯe�¾5D_��a,���7��h�̭��G9n�x�A
��c�,��ަA�
@7࠙�vy:=q��;�mu,ZN������'���-�+�U�J
���QC��x��9�a���u���:�3����m��O�Jݤ�AQ�����x��L82y0�F!����t�^��jۖ�8�{������*L�D�e���9mA%�w�P���[�&{h텹BN�n�(��ikՏ��G>(���:9�G��_ �m^kN�UNTt@A�6f�~�:�[���g�<b^����P"XuR�Q�&��r���k�Ta�O����Rl�ĊW);�L�Yֳi��/_t��!J�m�e�R��ȗ���%7����gQ�d�2�7��$>|~�3�jx_�t�����`�ݸ=b�=��,��g0��O}�����e�G��8	�I�-�"aq��ܿ�!Bh�lZ��4�2Dv�e|:-H[7���ƿ�c�l�d�\d��J��<���J}�����@�Kr��Ժ�>�����t�fIǿ���%���B���
����`G{�<C��R�u6t��1aѽ/�U��n� [~Sn7j�)A���a�2�7 HN��𳟪�,��D&8�5�8&��{��YY���89$���ȸ��)����W7ޭ#)�t�����26=?wY��z��^ї��Ĝ�L�C@�̣[��b��b��8=E��1?tt>
,T�|h&��]]�={�͟��!W�6��Y�prt��FS/��y�"�Z�ݟZ~ʧ�9�� ��y�]GwM%���5,�W?v������7!-a�.Fwu!���2�=`���nqY,����i�gl�]Lα���#�)ǥ���Z)�#<��O�\��!b���g�q���!P$AT���L��=C�m�;e� �@Z�����;DQ��15�;�#��Eog4)5m�I�6"w�Q�ԩV�q!h~���3�M��۾�1 ������_Bi�~(�P>Y��}����9$��lA��L����:4wk���)�"��@4��p_E��f��^O�B`�M���@gW�Մ�il��|��yá�D׹�P���_8��p�v4_=�b���_pg!qn�S��s�z��N��牖.��?,i �aR��5τB1��KԷ����(�����1#dJi�¡e�NS8{���a��^g����k�����(�d�G;��eK�r��b�^����1VO��1���c3�f����с�:6%� ��Oz���[ufJ���#+z�v�:bd�Az��	��Tp���M��ܔL��i�O�F���-X��"��3$��(x�h���!�	�ڠ��� ��R�%%Վ�$	�������N-���������ʭ/Ga�L��#kw�,�76�˰���f~�a;�u��������T����i��4��(����(p�i��Op�Q���6�ȑ���E��1�Es����V�ɍ��&���v�b�0�ȡm��ƈ��n�6JrS�GR��M<�?]8��ġl!1.�i^~/�����,I	v���ɺ_"��ǘ������F��*T!|���#&�	t���[o:�-��| E�;���j�}n�`�~�:��@G_�y�E�g�w��L11B��@k�J��>wF���})�� Vo�2��am��p���,p��<��3O*��5;�d��v��$١�N0�/��U�@@O^i��T�_ұ�'��v(W�c澄�����R?�_�E6����Ɋ�s��ۍ#�1�sj�������S������'�Fn��n2N*Ѕ�E�f��e��;/�Ն�V8p����g�{lT�N�x�^�S}$��N�������kFN 㧱&�j��%G�/�m���"h��/f)[�W�/�S٦���к���A�>G��pYI���FW����ٿx�r�����^�2(w�uf�/r�����y�<riw猽z��$��K̏)�8=�h;��g�Gh*��P0٭�;��<D�����qK��U�rH"o~�'�J��R����(�M��n��ŸU�b�R�[Έ�ф.I�@��m��'*�ʥK��=�U?\&��k�^�5��Ķ�1��`�ԬE�ו:�h@�|�� �.���G�ZZ���8r/F�����G��֦�8�k�#��sc�BR�	Ѥ:ž�ǟ%w�ũT�(����wR2��	*�P�?u+�
�\��b�^��$������y�}���/�ب��y��
�a��&u��GG�(��Ⱦ�3�⃫ɉ�ASX�cJ�h����Mu	R�b��k�j�א�gƭv	}��hH�����������v�춢9��CM�8��_!��na�u�O�ȝ�@"Kt5�Fr`�23�VT���r�e=�*�l7\�=���K�BEKk�tR����~:�	A��l¶<���
އB���;w�h�{�=��u�{�
s�4V���h �
��l�Eᖲ'�B�R����p)%�ۺ\3��t���+�������9�d�c/�|����o�dz9��ÿ��P�j߫V%QΠ#$3&�d���'pA�(ԁ�����GH�^��r��$��#o�5�n�C�R��i�rr�c�^���0�'�ONe�;
g�L�>�M5(�B�P0��șNSŨ��mq��4�J_�ѣ�-O�G��P���FԠ��s�qK���e"���Dw>ב�^~ܱ`Q�8��+2��X��
�9޽_r�ez�tv�0����!���u %yb�䖯�����`Eg�g�P�>>�B��J� $�C��W�;�!ң�R��N5QI9	׵YC0j���֋{��%�5��������x-&v��"�VΔ=)Q�y.�e��S��Y����Bvk3m>:����YM5�,��~��N3��V���Րi}�ǉ��7�M,QA�2���1�Gή��^���3?3���-j��X�r݌�C
>a���)�����OSM�p��f摔b�ՏN��h�:Vh�P���6|����X ��<�l�A���9tx0K�`��;)�ʇ�>���p�+�8�qc\�sV%�mb�� !dal�Sh��W,񣔬}=�2Hst1p�\�G_�H��[����ɃL��IN"�!�w͵5⸾9@��$�2�9�[w�{�����R.�[�!qC�w*0S�#yA�L�{�$^¡���-��'5��«�u�;�>�U��m �21���I����D|}�����22FU*��#>�6��������ᦜ̺H_Df�Ac���ո})�2E|�SU��$'gJ�헉bۯ�ׄu���/�1
�������$,��M}[�ʞ�HĀ&�I��dwI%+H��6GX�����s"��Wh��b�w���)�T��Ψˉ ��y���/�"����Y�m�����=������K�0c)r��-�ajy�(�֑�0@�(��~���lM�	��p��좉��<�h���t�� �(]��B[�9G&�����}HT#�Wٹ�b��7�#�����6xs����c+4|�k��������U���{��h�N�6��܈��bI����R��)k�\�8�����'
��b�դ�i��_�;b�r�(�� F���;�\xS�sAĒ�J��̀f���z���C���	0';m�f(h���M LT-Ǿ����F��t�hѳ�<K���E�,��G�a1��+��/��e���ʒ��Z�}3�[>�|��:h>&υ�`��je���dnjWJVx.�5�Ӓ�#Ә\9�����������
��[B��~}/qM�}��H�_(��_�� M��,X@3wB�Dy�N�� ��j����G��]�5�-E����Qfr$~:���Pl��քv��
%V����&�|�{'c_�^��������R&t�� �����VK���}"�����W*
>�U���d�p��L}��<6s�0�=��
�),-�w�|0�eߦ������(`����KdF��$���uo;-�*wA� tԓro�?X���N�#4��Q�t��gͶ�y���J�pS����5ǘ���JF���=��]�����d߹R5�.�(|��yr[^����$SK=�O}�!i��CG���Z=��+�[)�8���i�嫨{�H:v*t�I�އ?�h
i&��қ����v����!V-���^��ܡ���E�P�0J�1�~j�O� ���Г ���l����{n�mf�>��|S��h�V?���*{b��)l��u��� �`�m�#e�O2(a�38��Q��Έ�aL�j��Vt����5Q�����h"G@�"Ġ�d����ˌ�������>59{�%��l�3q��Ex��x	4R����z���*�噩LĢ�J!yl��C:�|z���zq���7, �Id��'�S#���xUyr��X��O-�@Vp��X��lgܡ2 �&`��r]\G�el���Hs�`W)��7�3$��(��ȭ��6���s�8�����o.��7��ME�cP�f�b	��q"kʎ�=_�dX��z 
�6��<�$N�5�ZA�J������~��E��w��Ϛ2��"c��:�lǇXw���!�岘dA��i�h���:%/803£�;��/dDTg���r<��,�t�LB�\t�R+d�DT�ƑGm����C`�}U �sYa���Ax˴."d��5�@�����qn)����	 [����[}��if/8J�����aK�f�F��,��ǯ��G�U��vǢ?p���@�C�>�9m�(BkU M��W����]2���� �Yh�4Sp������O=�U�'�/�������xt�$�q����b�w�b��w㬂�AW���8Z�^�������w��H��^��L�&��C��j>��`���v�Ob���A���/�`�����wu�Sn�ui���ZwO܇#���"c����t��!.��u�r��´�N�>NZT�j~_�;6��UT���ؿ],�툦~56n`�5���*�x�BM��Ba8��?ĺ]�\�_#�ѥ��mS�^��]�э�����Wk�bD�����5��'.��Bb��8B3���J&�0u�@�)�%�/�IG��:����U��	��d��ͽ�?�����Drh	�}�JY�{��=���:�Ú�û=�iV��\?rjo$6���kz�C~곟���1a��HoK�����<�S���P!/U� �/lpǹ�hb&Wql�QN�Q"gU�<��UTpe�YxĮ�ޞ��/[S�90�&I>���VAZم��8�?����\jg����C�hh��æ>,x�n�B�5�Wܳ<kf6��k�2*��������Pg܏�e>V��爕ccn����	_��I�j�=�7��~������m�����7��p��Q�`SO���:n<�O�#^?�\�`�s���^\j<ֵ�1�Z2h;�9��b�
��s�7d�*a�{�3 Xk��9le��h��	��V�p1����	ʓA��$}6��`��i���>ԷH�kKZK=�=�evl��*	�if}�0h2��k��Fjt������n�b���w��g�綛eޕr&���N2�>����;��z�B�Scg;����H�
�"N��z:5�)�9妯�I��F�b��?�Z�J�����c��(>�ms8U���`�����hU���n�5��$3��U)�x�,d1��衤�iK����^�[�Rz�npyܽ���d �S�#�b��z0��Q��0��5:��,Ǫ0~S�h�f��A`�s����3~��RRG8m���� d�S���:�g0:e�؞#�/�B�*�^0}�&����r�H��i��2�5M�P
#}��v��|)z�ʌ�]�e�) ��i�3򍉓"�{F�x�W�L4�8$�B�e�}�q7D ȐA�2��w;E�.��VJ���a��qkaWy}s��/��#�#0T�|ψT�߻A���Љ�Q��@؆y�Rq ��ά��������-�cY�	�x]��7R����q�nx�0�)�v+���*��-���B5�xc�o���:r��A�n�d��X��O�7( nʥ�.���Ș�X��6|2��y:EQ��8ګ�M�_�m�<��=��[c�Bwc'}��Kf��e4.o�b�Oq�ݠ�(�`��� X�����G�s3� 	���3}��X�n~Ż��r�m��4u�Z����d�VA�҉Cn��'�j���y�t#��4|��3���TCJ{u���u9�x�s~�����(�t�};�X�r�ڠ���W#��4�ʠ(Y��1��$�H�.�$��!�??u����ڣ���4d+�p���Q3����z[���ģ~���/�cg�.{B3�G�ַ���=�Y�sS����\D\�j(���f�$%�;�a�hl:����DD�K"�8��z˵svVpo�B[X��͍�L��$x��۳u��}A���� ��<Z�;�ڇۛ�ZO�������d�7ԦU�Hw������_��욁��^��ө����N�:����\W���q�3��b����<Mf_��}^��)E;�f����uCXB�S���W�8y��+I(�/e�1(L�A�+I@��!�gl�JiZ/K��sw!���! 4�ӏ�+��b�����1�g���V�%�vsĞz��-�kDw�����@�Nț�q[�-徆��Spy:D�
8"|C��
ˆk����=5�!z[�!�Gh�k`�t���!���o"��2U�s��
����)�y{�N�2 ����0E�[;0�*���:��Ɓ�)�+�f�J��U�P`�J�濜ޱ��`ގe�{�U�#}��|-"�(T� ���q��Y�D	}��6��Z/��O��7U��XN��ܪ&�d�t��>Sř���8۠�X�"N�p˪�Tj�ؓd�2(��g�F#�<s�1�]v�N�I��H�h�e�ܲ�$93E�HA�§�ړ*�y��nntbŨ�(�M���<����o��CC��DoaΙ̰U�%�~A�츉�:�-^h3���t�rv�i4����3� �Lxi���e�\���p�-n ��\���������jo��Dm~(^;1ӽ<bKU�~��/#�|޸��qW�8��2`��[,�+r��{����/c�/v��&����B�#�s6������i�A�"($?��{ܫ���Δ��c.š����xWB��h^��\��ڎ��0�̏��b#'�s=kͫa��#��^���0�Ը�=��3���?ڗ�ڿ��51ޯ���^t���YP"�~Q��m�*;��Zd������W gܞ`�"]��fn�[Y�����H��&������3q��r�'BT���C�p2{�S
z�ʦ��7�qRS���<�������J���� #J�u�bS��D؃�ሰ�ڊp�&�f^�����<M���{�gz��kଘ.���X��CRֈ�i�lL�s'V}��W4��@�r&�~$�;��M��� 3L;���~:�Nc�cϷO�dC��eBM]f>��F��Fә�_릋H;
|mz�"ZF��&�y'k%���=S�.�5n��nX
�+�4��Lx}�n��Ed�$���FFH���>����.�uj��}1�}�#e������w�8�'+�W�wL�C���V˛�qW�~��jW�|�ɳ�dnN ʳ�+I�
?�1�'8͵]�+�,���tۋ��$�{��S�V���sC6
��^s!	��;���Yܱ���8��ܶ�o��q�|~��5�5�7��]��Wl4]��MM�H$����i�$x�{�A�;Mu�=$?U�!$�ҝy��TD�FܾF�͵��V�r/ݨ!0zo�,<�Q�`��s�� �������c�����,��e���+%4ݸ���ıD�%�!��jDk��;��κ�4�T����eq�A�����5�~����W��1�W���S�FY���2�`U��3�s.�ܩV�P�P��>�B��Ũ�z�l�^��RA[zFN=�L	6B�,��JR��WQ�<�:ß��}�Ѐ�ǑV�!��*���O�CL�oG�H�Hk�A
 �ʛL��߳Sߠ�f�Ly��=�3�(��l���b��t�����K!�\3�iN�~��&ѻ)T��p=7ˑ�r<�˧��~�\��>���bt�_V���]�A����iu��&�_u�/��ɥ��rϷo�\�t�{|����#�3�ѵ�p�q���C(�������H+�L�,��$\�P���a�
9���\�k��������W�Rhr��ˡ����W�l�6��c�ټY�.�TY���ӯj!�t;R���F���r3�d��`��� �`�&ʻ�x��-�����镇S�ۦ�����Hv�c!W��@��!w�%u����J��JE7o�$���O���e�J���&#�C"�M4-�~�m1Ea�&V1�ūl�b6�y�G���C���&��41�_;�!��7d�~~C�ƌ��T�L؆�"��ypQA9�H���30Y3�������^
Ƌ.���
���V�ñ�`�6!ヨ93Q��"+Z=1LX���"�����2s��,���W3H׆�89�w��j���sW�v�mK��"Qei}�\]c�5�D�r���o��!v�����7\�;ly����.��g�Z����������Р�YI�?�׶��?�W/��G���=o%&!�΂s�[� �HvMpVTNa����N��.����(�i��ڹ;�7%��`W�Qn��;#�F�'�t��`�j�O�]֟�>s�ln~#�fu�q���h?yC@lK�Q[���������{~8 ��Id����Xk��' ��~V��b3Ih�0r#��ɫ�hziP�#��v�(d�]оYƨ���"�A<�U2T"*p�0�9�f[doR".qjR]����%b<
D�X8�̹`�:���o���D a�]�
gxgg��8�/Wғ����R�\�ܞ"���:��pb0#��uu�h��4
����|I�N0�L*X��&e��S_�_еíez��nyq�Cc�a��,x�~�c��w$�oD� �>��Ԑ���CW�p�X�3�R��S�U���wވ���\��zQ��er���n��
-�p=^��	K����/��*e��\i��.Ѩ$�.PMB)��P�U) <&��/�(������2!C'd�[Gl����3$�[g��3�����������5yd�V��hI�����S���yn�`�n�Un��̥LʄKQQ��&`\�c�6�;��hV,��J��g9x/���x�8@y%�Wռ�ƣ�a�$��B�l�A��y(�|�H��A�,]kˡ�B64�7p����3q�I�[=�8�`q���v�ׅ��Bd⟗� dq�ƒU�d9��*�6|����6&B��C��13����st��vA�{�R�}�� �S�X��9:�/Y4�O���0g1��Bd2��.eU�GG�)�N���x�\��m���8:\bj���C=�6 ����w�h�;��0��]��� ���7\Pv�kΔ{�Y #�T�H�V��V*}?�|���I�M����.:c���|�_Yr�u��B6�~���΢9SL�>��-�[4���� �Ӛ���%9��� G�(�������T�����R�/U�#*��0?l�^�յr/�g6>(��g�0��J���� cKXf<"`���ԡ@~�I�cų5�:�\�]��G�t�����*A�y�� �Fr���¨R~[�f0�Ҭ�#
����'�U��"��ti=B;T�d^��ё~��p1�Q���~�B�C�!쩗L�Aͤ���c@�������a�0*q ������
�Spl��t��D��!~��V��s�[�Ű.��2l,�&aLk#&u×�c��8H5v�X��:._}7]+r2���!�@�+1Av�{��҉�h�G���
��
B�iRc���$d��/��v?$���6�(�O�ؒ=N��M��N�1�kvZo�V���h\�m��.ޤ�Tش{��>:�Өg]c�@JCB��G>s��B�ǛX��������Mg���DR�J������z�}Uq�Uɋ2�l迣\?wD���ů.^y�8��4�~�.��/����y;<���7~2h��2�. �w��0�`�,4��ۭ+8�o��1���H�i�8�A����7"��U��������-c����̩�/�"����&�r u|S�����f�p|��G�,X٢c�b�-�l-��� Y�{�Y�@/]p5TI i�wl����{��`����9QT+)ܩ��%9�6�1�,�QS�/��r���k�cK������>�|��$-��aR�ky�^4���7~����c�p�n7׋�+�,�9Խ�i�_/���D��<h�Ƿ���<��$�틡<�0:1��hg`�:�i-*�}�*��ͧlKp)L,�%�Lf=Z��1*�#jzB �ua'��s�"L�������~[3rM�y�ۈ�q�a��<c�H$� �r 6D�� s>K�?}�s�O>y�E8��wࢄ���<�.Ƴ��[�m�~�!$��Sr��q�'����N�DƆ��I�@�#��Q����E��])A �οτ�~Kݰ�F����r3
�Ǖ3�H��]f�ݵ��	������#�a9�>z-�-�ĕ�D ώ�uw���h�W���>oF4�)�3 ��ҹK�(���/�}':#�����'��h�ΒQn���U�pVt�̯b���X�إ�eҩ�y��ڜ|��C�5*7�	cH�e�&��n�ۈYQ�b�~�V�1��|����q�bHT�>�J�*����J�ӼK��-�Vn�Ԫ��iv�ٺ�bl�������o}q"���>��W#��;�V�%J7�ް'�r ~�X�\;}���z���"L��]%E���:l�I+����t*>d-Pp��0���3���7��6�5�1vh���6Т4!��X�by��a�׾�nb5�T뚀��.�~��؏�;��<˭�L`�	�GL�S<�=�tLb>��wO ǸZ����$�H�{ߐ�`zi���<)5��<��,������!V����D;�c$@~��*�f�����&�B�T��S�Gd.UD�Z��qT3�7~N��L(��U�O���.���$\�1-����g���  <(��#&o�N�GR?�ߟ�ZܴY�sz'�L�=_k�r`��$q�k�|J.�=u��f?G���-���������UY��Lal�	Pt¬�yo�h����)��vm�o�p�pZN�̦6
p[�f�y��H5p���N6�����vKˢ}b��6K5�Ü�8ߺ��R������a��Y����m��r�b��8��n��y)'hče|�F�,�o�� ����>s[��T��|I��X�$v-�Zd���Mqr� ���Y$gԩ�sC]�\���e���}7i&�����/�.�_�K���H�㨪1�K�ñHk���7�z\j�{���"��/�_v0���5P��NN�-$��:r��Q��\Ψ:N��a
S1� �>��ܶ V�I�A�SE;u~�Q'��\?
�Vi\�9��6�%a�"�x��&{_��$S$��m]g����ٴ�X����z|k��<�Jr����Űr��PK%ư�f�ײײo�h]��������	7���9l�Mz�0����,�o������Y�ƹn���[:�Bdg��#�#D"�t�Ah����ļB�Hq�@qn>�ƿ���4$l%:W\��j�U~��E6RI��n~q�l�42�ųx�h��ᇼJ�+�ڡ��ʌnl���U� ����Nܹ�QkX�	�k�"'o�bp�j�m�]|V,=:D��L���L-o�����ju���+3�8� �8�[31R�J���P���
Q��KZ|�l�:sP��ժ6}ԬU�9^G]�1M��\��ߖ9���t�ϖ��
Gg�P`0�yI�bæ>�&3E��3u��F@�z�J����.�6jQn�@8>AoECF=M��@?�dx�拽��@�K	���.3�ܐ~�zr����gS��{��5��5f�;:s�\�G�M�J��!�ʪ��\��W^�`����dn�P�s��qi �Hdzax��W�=^��j���4�b��M�y}����61đޖy�z�Cac=;�(_�ʻV}܃��+V9tK��n�ґ�������ǖ����e�3�����v�f�\SuЪ<?0�t�m9R��t!z�~��i��]3>
�Dv��[Ro1�bj!�ӘMS^�ωk���!.p�6ߑ�T=Ls���~@����$�L�φ���+��6��pD�� ��r)�V6I	�*@��쇽:��+���
N
���Irz��B��p]�TOȎ�4��^_U��y#tE�TN��~RD�4&�ʜ��\y�����K;#)�ĥx:Ɋē�k��9��g�n���0�u��\�e�фw�b�����k������D;�A�U�66���.W���ڸ &�۷�#Z����~�K�q�|���rWv#ϩ�r�fm����1�yX�u�n�Ng�R+넻�3 M7��V��h7~�F�؁�Z���Id�����*�U<���C��>CNn���#U�ک7ݠOB�9I�*�l|�rсU��9�
9�m��fsf{���G�u~��0�:3E!X $�������*[&5�_�6��r��@a����T=���k� ����WV���K��:|N�Xw /t���5���3V*ޞ��P���̄�+�^r���}�>�DH��ٰ�ڝ���H��Q����E��ok#��A؀�<��I�=�I� ���b=�Zq����J�w�g��Hm�=zF[zgi�Ɖ}]qާ"kwMp�NG�����[��_iXƭ_�L�	��r�����j�+����r�dը�����ז���"j�MO�L�,�p����
וj��72_e^���=�yFң����yT�W�1��u�V��u�g}�((�ؼ�2�g�O�D��d��6�Ȑ^ �Wy~��Ǘ�pe�9��2��#���ϻn�S��V��.xBc�d�i����.�8�	�������Fx�_w������f�в�`�u*"9+���X |�;�8B}���
��!W4�5N��L�:�"���']����aK��MX�j��ؘ�M����קw�:��}5W�M�Am�O�&�vW�>�a �3Xe�u_�g�)P.`��[�!��20��2~|�_-� ��'�޳�yVe�/,�D^AZo��>+��}�]҄���J�-��f�p��1�bF1�j8-��O�KK���n���3:/ $X?�Q�����AcF?cLb�09-�=�y�2�* L�r&|�܏\^�F��};e�"����FD],��|_i��í��/�rʜā�h�,V㙎��{���ZJ�F� !E% �;2Ċ3����n�D[�<HӆX���杈�^�e�Y�BPL&s��iQahT�y��k�SW�=� �����>����%3k�O�L�
/�ޖ<k���~�Ӻ�x����Ų�?IZ��e�Qb#�_)Qj�F8u�| }���u�m5�<yE�,"Ƀ� �5�&�zJ��nS�w��#�`25�<u��ZT��ꩣ>]8�y$e�/%=k��#��4����髩�2��!������q������F��V�W�-�z���s���
Y��Wڴ�/U�P�O�q�W,�\[X ����j�$pj�0�J��ډ�CWz�|���0wd���ҋ�Y#�l@#���wN \η�ٲ�x��:{ۖs�<Dv�#�v	����oQU���5�KZ1ԓ�GU����N��1�L��cBQ�E��'���3+��]����bKb1�'�ާ8�8V[:[��E�EIӌı6m��}_����9�D���h	ғG$$ {��pg�����>�<�ͰU�#@Պf����Y�j����>�3����W�Mq*�W�32W͇|�@��%��7UH"����'�2�&%O�޼B�1Owc��,!�5�%.�d%���戈M�!Y�����o�F@�;Ԩ.,>	�y��[4r��!d(��^8��"@9Q�x�N��ر�0h���W���k T��ĸ��T��E���\���R?�lvf*{��'����z���%��sF�G�QD�w���J!ܜ5�!��k1��0�~1��}�S5gģ���G�FZ���������C��'H�
�7OUnGU)!�� Gٚm���R��댃'�m~�Av�4t�}��q����ngݞa��1X�GHQ|�d�iU#C0�kr��ֻ�sP�� 1Zչ�E�u����V6�����H�� \��^H��~���ۜv�6e-551�(�c8�ptP_��D']7v�}���V��d[v��<�E=H����m���Z���g���	�,tؚ���t��&���>0y��&3�ff�,�����(#��>/�Ds�|P$��=��xߐ���"%h�mCcĸ7���ܘ�/Dx@�]U��UBT�c���q+��ܒIL�����o?pN7�=gRw����h�t�Da���W]&��=��X>c1W};6ϓ�M�i���QO�cT���=�����Ș~
�p�H��<�ř� k�+ \�?ӻ��/p,�,3��|j?<�@�"��0Y�>T��9��^>iت���xF�D}j�^�R�Ɯ��BZ�m��C�W[z��k{�|����̾^��������la��g��H��U�f�>�t�_��A�4��Vm�Tvc�����|���j;M_T��,\�gq*��֞"GìL<�Q�B�&��)�c/�ѡS���o6j%w�~���	d�9+t�A �����S��N%8�@��lƞ�%����k�a#k}%uv���*�r��*:�Onp�cᯠ,�5����NX��3�;��~�Դ���/f�ل�*�ڣ�qMՄ�l|�K!!�
C�cm��M�pe�E��%�߃`��xoE�����^�{�x@킠�g������In`s�0���l��bD��m�An!M�.�R�r��o�0��� L���w;�L.��%j�2�CK
�D���cߢ�pРT�r��BbI�M�ـqŻF�K����_��/>M�$.xg�/@f8a�2����W�8ŌM�[�3^����GsE�/oc�%���.���@_	.;�ν~P�"�@��jrDW�! �m�/nІԾJy��^�zM\�s�|���x���h��G;��(�f�� cA�����&��a�IO��{b���+�����=�r��߭���Ɣ"a��ȉ�Cl�dޢ�y��f}O\G��^�k��۬�]�3�`��:SA�o7��ͪ}���+�֢�}��AD9�É*@�]��P:�4��6�R8�e���
e���|~/�9r������5LÚ�o�Xh:�����w8�#/��^����	Y�V�l:8�vʛ�E�U
�����?�[��S,�o+ ZϘ���&%�%����0C�N��M,��W�U���\�=��`@�����m%�	3Ƨ
zD+.�n�Hx�����8�9͜?�r�W��_�n.�
Ä�<�˱�;��a�i���T��Đ�es��o�&�xXn~�*,~,p��+sj�7ZG������M2<���"*�qc�m7m1ĸ<���е+����&�=|}�����Lr�Q+� C ������I(��\�Bk��Ҡ�[r�T#�]��C9��>����&Բ�"�Ut`$B"̷��9x/��6@�&��E!��>����������u.�W�Yx���lo�������Z���f*��{��}XrMW�L����g>���쟑y/����őw%���~�аJ�q�f,�Z�.ˬ3Y�����~a��1�}������,MT��Ze�s�8P&o�浉�InOK����kTP��V�>������0vSCæ�>�%��S�%���,,:Á���<����!j�
���f���� _|���V灇�>��Z��Rc�G���O���\���� �8���p��!+������P�Rѕnq��^�T���\�:M���Ķd��|H|�38>��s�2G����	�%P�o�Id2�j̦��NB~����z��/�)�u.���J���aL|��fO�u�-�2�D���>���y�<��3[�'Y��q,���$��a
�������p�YB�+��`� �F�!ߣ�� IE��F'P(܎��e��ߨHM�M���e��Z��癟ny�����s5=1��m8iY�Hv,r;��6>��\�o(m��-8b{���k��,jXЛc�|x)d��3�����+��y��.�B�qֱS�P&�?d�Iy�Ҽ��_F��zH�RO@��K7�Nb��
��E�S:S�����ʯu�r�)	�G�4`�����g�\؎MSI�w��{��c�L��X (e�`���n������f+LǦ}�X8�t���(��֙|��7��%ICp�\32Ð:ݗo+Gt`D�5(fL� c��s�WR')zo�y��+h8H;h�iAa�l����dB��ll�u2���/(7M�٬����A��`�e�G��~GÅ�3��h��b�F�VhR�1���b�y�դ�$�3���prG3�^��}���A��/�`i���)۾3A��o�S\$Ys�]� R+h%I(T�V@#�� �RO'���"��-����<��8%sR�	P+�!�Ѻ��#�Q< @V>�خ2�?��6j#������Nº�?r�]��O��=�p?���>om���@�s��Ꚏ�����vB$ݺ�7�b^צ�m&�����x�f�U��r �)�Q��J,Eiˆ�ͭ�=����!����&s�\��6�.M���*� ��ژ��/fmR���!?~�z��հ���[�<��.�㲁�:���͇�_��u6�D����P&�JaaG��c��5L*=�
m
�[2��.K^Y��[<f@�����+�?;���Ez�z �@�Ŀ�WS�uF}�U'{#A�y�*��%��dx�nup 8�f��C0!�kZ�I�o��_rTs0��` |n���  :��b$�H�s��T��*�v"wnG[N��ņ\�q��|ѳ:	9�E.P�����'�lS���@aAT%E��n~��~Ղ�F)��j#%|���J��4B�`�y� -��h���77�m42Eu^��S�$��4wݒ:�G�OE���*h��-�/���ή�8!��Y6�\"A�NG?ڮ��~��iB�qL&1qR�Ԯ�
}���!3�Q�q���hM�\֯�`�\v�~��Ŝj�'���d�M��HRl!�t�ݧ�p�6
�Y�HOv�za���~[� ڎ=DR08�_q���Vh���.�a�'/�Sȩ��v���!/���z�e`�V���[5��W�*��
,#t>����<�`��e�w�Ȍ@����Uc�|Z\������'��=?>
x��#6{_X���~�-�ł�[0������U�~7;��Y5	�}�O�F׬B4-�_�Q(7]GJW)��uP{#푷��$"��l��8lwuv��BbZR��x>�z�?���Df@� ��	�2+���:n��*n^�A��6~�8kdӢ#5$��/S�L�`SWQ&#H����\��Մ��ú�=�A��\sO��f�S!�`�k�A���YO�M`T¼�@�Jp�����-w7 �!-��&7~-�~��E8w�@d�{t�V�ԕ�y��B���X�a������Q���DPQY����q9�Al�wgLoK�܌c��IG�C ��8&��(k��"��_\H�xo��`�J�*���7=�-���2� �:�|�d�-]��`+��9+�ͅ?>�qj�Jք�|�OX%�P��Eٙ��a��#��<bF���׮�*��q.#q$��|�v����a_�~�C��cl�L	�&��rj����j�Q@�IjB�
���ƺ�����#k�/n閨��i ��D,��D#�W�_S�c������?1����h�Np.S�=��p����͏~׉6Q����Z�71�Q�e�/gE�_�~A�Pu���K
�O�@˲2+���|��v�id���{�iozV@������J��ŋ�������,]Mw�� lsB�[3KإSf�z���h�/©�K����#���oZ��q�Qd8`�`����z+Y�Y�u����Oq�2y�v��,����X�c1�N� q�J�R<����P*��m�.���ު���%"�q�B:�9���C;2�[p@��&��\g���_`��Od�r��;$�@�IJ���ڝ�܉lo����ݔ@	x�E��hi��H(�otube��e��
�à�ݡ'��[�ȭ�H�u�A�H�Ѽ�����B�#�+�jل	�:`ҿ^!�.RE�7�릍7:�}Y���sR�itU���m@m�̎��[g��+����~������c�D�5/�ݝa��f�1%r��f���.����6 �J:��ѻ��|������[,Ӧz��4��@Gزwa�ץ`	��L�MU���5�»�(ώ�U)��]w�k��Ln'�:�!o�������hC�2��+U8���"�W�ǜ7�# �!^V �{�h�D]�~>��M�Z�P��%�!gV���4�c�jE8����?σ��>!��|f����>1��u�P�]<����6�,kF��G�)���L�n��(��0ݢ����Q�kj��Ff&�(͟�W����+��Ulo((���3���R�-��������8�	i��Ǟ�Qc$H�����14�\4�)���9���.md�P��O������D�o��ң���
��'�*O�ӎv��ztt���p_�(I�����R@��YaK�AY�#��l}��x�Y����u˼�ƍFru���h��.�ͤ������>�l�e�oq���B�V�aF���u�,����@��s����s�ɰ�J�Dd�!�Qx]���8���p�+<CΕ�<�`^6T�*���T�e���R��:Ѭ�򘥳'S- 4kG�݊��>�� �w�U@H���SV�)�OC�흴�[j�K\б�b8�����lo��e����t(W���j��A�x�-*Jç�"ۓϫ^Ӌ!z��[��V����ҋ���s�F�����U|r3n�`�i�s��cd�)e�-9؆�r����ң@}���!3քЂԥ�rp��Om�L��y����R��h��j�k�Р*8<i�U��d6��}�8@<h3[���u����q�1��zK<G�����霜�ׂg�2�dZת�W-3�e��.Qĸi8���ZuN"I���kc<6�� N�>��e�����RM��U�4�aѹ�,�����fPCKO��&c,4�������������s��yX�jڰ��ڈ�	`�-�L��5��	�Z��?m�C�a�S���3V�����7Xù<�q��FV�_Q���^��zij����SW��/sS�t��	�PW�3���n����ޕ�q�uU��KH��>���*sO��Nm�5ȃ�@�����a��PzJ�p߿2���>���4B�׬�x(I�l:E���,�PPA����۝�T���j��mdK�����()L^>�Af`-&yY������|�w��@�f�H<f)�_´LO�)���N�u7*xs���é��X�B�+�QP?����g�>���C̫��(u������ÆK�A���r���6_k��گ���O\Hb�Uk����=l���������Ĉ��s��m�e�˨d�FkjR���G<t������_���rz<{�% �՘�=��!����}HLj��l����_�dbV��:;��Li�uκ�+�,�0���\3y�%�O������͆oP����~�����-R�Q���XǊݤ��Q��/Y��%�-�� �n�`���=Q�O��[�*�~�cu곝D�gl�>e����~�E����]>|P3T�p	<y��N�5.ܓ�r�u���@ަ-��[�
U��a7F�}�!8" �D�D��	=Z�&W�e���}�xk$�3�~��$aӭ�Tً\gTM>�/E��z�xY0D�1R�����Y�߅��U��ͽ�C��.f<g���)V�W�R�cc�	�h�м/S�� �&YOrr���X���%��|�~ 1��(}6���fC�.����b�B�NX�)8�b��D=�$]֪6�/a�r��2�=� �ba�B��E�9
���9���XN���J��q�~a 0�tCAoy���NGB%�	r���
lg�D-9��MV�6j�,��Ѭ��uz7�`������#�M��ж��wV6p���G4�+gbVj�
YRF��FE��c}/rDR��﹆�߅w����]pBD��4��tGE�U��G�n�=&���"�e�
�Ч���o0ӏ��#?��n��D���i�f��Q�r(F�������<�0��u���E������E�#���Pq���m�哾���J`�B�i�
nc�(8��C��h02�fZv�g<U�X�{Y�F{����y@��SP@�R5?�	�R���4�o��H��Y��2:@�#�g=%x�Y�G���,���v�ljP��(�yY��=7Yڠ��G<՜��8�+�~4����ި�Fr�s���&nν��B�����"����?@�'u�ذo������~px���!�����}UsMEeλq���!��\!�q���2���*n	�b?�/�E���W}#��Ǯ9�%�`	@J�d��n���/۟�����|�O�Rݙa�y�Xg�Ȓr��ʩ�&nkziε$]Ǚ&�9����(��H�ᑍv��%�9�
 s>s�NX��xQSU.,�ݝ�R�����l�T"�r�=��A�0ƇȪ.֒�\P���9.8�C@�;��6f�#�#�e�8�=��r�::$`��� ;� �zi����f�n������Q�@�!�6��E��V[s�شv>��x�B����ф�>�a9sc��3���A�\�sAj4�i�.,IYi�
�C��\��.l�]�U��F��8��(0�J��+0F%|�f�����~����q�6)�l�1��@C=�:��{ȧd���\]p�ݐK��2/�N�}��#��V�}���>3��ܝ}WJ�R>^{>�7�|����!+Y���7��m'������[��K���vK �E��W5'�����_�pŮe����f2���};����A8��5c�޻^%���7��_N=�a��(����u-Y������>�A�4�����c�����@c��4#���<�,��x��2%���BϮ���x������9wl�	����0!f���g�9��Ðc��ʇUPf��n�����#����A�W��!��)a���۶�X	/.��^��*�᩹�m-�V��g��O�7�T��9���XoYy��w��ťS{��i���% �_&�;zm�)���T����g�5_���M���9�c-2�8�˧�K�Te ��h��	�ˇ�z�m�z��2PO�lâ��DQ�"2b!;�v��҂�&r���d���1��"�Y�?J���<�ĝΕR��x'�-� �V ׌C�W�&F���-�&���_�Q3x�T�����������x3\?�},{W ^������۵�ƻ�sϓV�&�
�9�\� ��K����E��q`�շ
 Rr��^�Ԁ�N��}��	�;4�ֵ�fp�؎￰ύ���36���f(��GCx�|'���������h�7��$���L8�����B�>~J�j[�t���3���&�`6̲>7 b0 �s!��ϟ�,�Tcy�@*�TJ���
]�N;���[�jDH�`� w�l��L�.#e׳�}s#�B��3eD5� 0�����B\�~>��_�)�S�77��y��w�'�$i�(����%��3FP\�z���I�:Rx}��a�Vgc؆����9��PGY�Wa�/!@��i} 1uS�U�7�T�r�b�U�G�,�".�}��x�\T��+@�D��gy]Jx�^�v��JK�c.!a^�)����@~��`��hZk���3,��kZ\���}����S��=t���7����Y}LV��V��%"x�Uq+)oʈH6�[�K��l��s)��5Y�3�����)� ����sX0,�#�{�GB��WDnKP��-6Ü�i�[���jSd�ȧ���_K?>�	:��"��5Y���[���<LA3 m��˚!�F�߬iMH���$-�e[ì��]�8�A4V:�k�oJ��h��)������c�B@�1���Ƽp<�r��Ϗ�	�k�I�5Z�ج�G�|)RlE�������],�������?^�*0�&0C#;p�쬓�[���V�p��=kي$7 ܻqa6������6L����$8F*A�lM���񩶉��r� �jM�c����U��]��33�P����P�z}3��x�ٰ�;lJP虓��t/��Mh��%`7�Ϻ�Խ��/z	�}X�KMf��|�-�yg�GՐ�� '�1�hq�H��ӀjJr�*P��Z�+���ܨ�u[��
��6�d�������"À�E鮗?����;�m�#%�|�*'5et�5k	]�&��q���L�'o[�iB�ET����-$F�E�� j��������=��PwMqJU�;��?N���@~�ħb��n3��Ѯ�Y;�:�Zl<* ǹ���e�`�v�j�ay+�0�Y�TUς%Z
q��c���p��F���3k�y-��,�
I�KM��)����»�C�	ٿTզ߿�2n�HH�����}�]�,0��/�Ą�P�u�<T΃4t�IOy�������R+�^�����@��>�f*�),�Ø),�M��ӹ֨#X8	�3�+����q�n��&�tY,c1!y\�w��#~������ڤ=�l�(��.�������D�O���Ŝ.���0�bha�wn=��B���F����Fʱ�adp���{ViyBt%-e�o���M׻�M�D���4KݮR��l��#"�r�����0�B�[�����!�ۿ�@'��q��\m}FG2�ؚ�Oʐe��P�-��5y�"������Z�J�ZAQU�Kt�M��4�vu6v��g��BɩY�w�Ǵ�=�j���ڽC�T�����)s@���;D��L���_���U
�{� ����jA�M�u�`kgI�
��p��U�3�2mp�n(�y'
@8��G\�W�\`��w���9��V��(��N]܃Ńx�1iu�h�W���Mc�% ����͙�g=��,�se^~�	�����I��_�)\-M�	�x���o�/5v���kT/�n4Y��$��j߃$������Qm��;�<̎�����mM���AM򳬾O�ͿŅ\: o���i�~���g����u���E%���׋a�]���
ra^�aK�X�J?���X��zEF1:bZ�[NV
@�_�q#mP��oEUA�h򈡡�)���o���޹�iz�1������1��^~��L�����g��b�Ӯ��|�yWc�n]wuI��|��`:���\i���,�� �\�8){np�y	.AJ�<�$�5�^"X�nA[�K2�
��G�vD�r4jlD���rʠ�{Z^Aj�?Z4�f����T�_�ɓdu=�l֛�
�פ������A��.�S�>EOn�����5�M�It���I)����,�3:#3��*�ɠe5�@�j�7TF���% +��Ĳ� �T���s��b:�	6h������%�3m�4wb�@T�@�� ���iABɽ��`��ë��..��P@e�ЖI��f��e�Tn>>%.s�sD�����F�"}g��J�E���˜c3�U���n��w2�ן�w:�g��~Mb�0�l:*jt�j��K-3"(������k �$�'�A-m'�=gPM��Nz'}��i�_�AEN��7����oi)�����W<��c�ΫG5;�Z���n��9�JS?��W�
�	Cq�02-�q�@ V*є&�M����l����i�eϵ�BP�ĐA�.a6 �'71��Q.p��-�q7�E�5 �������Ό���9�o��Ih�� dAY�E0���a��YR{���C,�%�7KK�IQ�II��Ed�^������Zi���`�z���%�#��rxJI��f�Ĵ]Ba�Ѧr#�5�H��۰Z�-���%�b/^p5m����
�q�M�K��o�q/�x-�`q�*�D1��&�>[	�K��B�~�G!/ִ�?�c�a�*m�7*�SVv����IƁ+�q��F~�eR�"�hk�;G��Ӟl��*��Zέr
�I�>��C��XP�{���h����B��� T��S��p'g�B�C�0����W�7\�ǩ������i�rM���٘٨����~rC�*��;'/<l�������m� �N�'/$X[֯����;��L���e��v�ؖz�E�	��6�t�w���%�9�Y'�R�jSp�����%hQ�﷓U��ԓ�G7�́�=��/��7*�d�ڙΪ��}O�nv:q���X�T�џNN @��{@e$Aқ}�2��3.Sn�dм1 di6]��B-����&�𮚙Lz0_qg3�"�<6��z]j/_��g�����7l�nD�]�}���@j��Yсf�j�T:d4�s !CH�G�]����Q�Y��Q
��x���
��C�X#������4b\�����o��>�̲�Q��V���-Q���lR��&�
Ro���K���F\��g;{�<��Nm|�*�Ζ�t��<SW�
z[�-��qc$�7��6�6�l�P~M�x`���C��/D�Ή��CZ,P��������j���� ��0�]��>���˂S;�@Y�X�2y:i `�nf�{�"}�^Zɓ,G�kɑFf�A ��3�a��h�z�{���57!�>z�M|!&�i�Ag N� D\K�$PR�=�� �x�4��\��N��Q���@���v3��Ԝ;8>w�L'x�9^�l�$ĕm��f.r� �쯽q�GI3]@ �%hŃhLO��X��}f�+��'����Ɣ\�&�I��R��xw���3�rܥ^ҷex��%|�w:�%vVrc�����ɉ�C�B��٧R�sIGwJ��3m�:JEU䜡��Oǅ�7�5 �tO2���K��9i	��ٲ��<`�4��wZ�ZE+�]�����3��T~����'{�Rދb4~��f�L�������i���j�t[tZ`�cԳ��U�τ����E;c�K�*}	��F�K�X��q�=����:��k�n��I<���[X\*�Kr����)����-��@
���$>�fuRbp��l�ҊG��O]�ܬu�l�
c��/Ÿ<������v�~g�uK�k<�|&������_I���d�	�`���wԾpJ+)��̚��b�����aP��=�M�|2@��|ğ��Ѳ��0�s���J/��K���횪�e=�a�W=����=d	MS'8�r*\N�T���d��&�
������Sp$y����:���U��lM-�S�)W��#Ӽ$��1�P�y*L#�����;��(VA�2�=�sQ��, ��C�W�o�j�&��g��Y��p�J}��{���$?�LN�'h�!]&5�����}d���Ye��{�"+�! (s1���Qwk� l����PI�c=�&*�_8�YD�0�MQҏ҃>�G�����QX^Yt�19s9�;Y���p����T7#/�����޽/��!��K�\��n񵗱~���V�	����P�a�* 7�|��U�"���c�L�;8-PO�E*�����+�<v?�̌Q�V��~�!(^��/�(�I�������������4��vҋ����*��].
Ɵuy)T�5
b�V��m���[�=����?";�CIFܡI�%�z�/d��8��,Ѿ\����W��]Kē4��+�4��rγ04@����J��	���QO�ڭp�+�1L�O�}��.vՉx�md���Z,Q�k�|LfK��L��Q�hIJ�-��20�N;���hV�GEk%���>а�6c��ɧ�zLwdR<d�!gno��+z��z�����̹�NAn)�Ӂ���~�j:�����v$�Q	�B�����M��*@+Z����7��x����J'8�6Q���ѯ����yː�D�A�2T۶�\�t�<[�x𛥅�PoN�L夁�(Δ��|��Z��:wX��&Г�!����NΤ�UF񬅈]�!9q�#�6Eǿ�R�-�R���3Y׉@H!	o1l�T�-y@mL}�u+eHMK����J�5�����.��S���M�'��ƪ�<,�N,/cb�;�&ZNJ_ssEq���t�����F�y��YY~�/l&��P2.�*�&o",���V�FW�V*��MH�B/;�b&�}���S���	�Ȯ��[ʩ��?����!�#����
�ͺG�̗�Q0�ԃ  ��6��H� ��p��<�2C�Tz�3)hn,ܟu�|��8��ְ��Ă���m���^��)+��F�2�j�joN�ҹ2�	Fs��F��ڎ�y�	&���piǇ�U*�k|/��d��A�<M��z;�]�Ec�,���)���Ia���u;��4{�BE�=�&�Z��4,�!����O �<�B���ȇD.T ޯTB�/*�;�Tk�SM`C���d�,��ڃ�q��ƭ�lw��j˯�hNh��ο�L�D���C�驤�eM�ìPN����U�΅�9���y��Zc��]F�N)�{/rMz7����e��de�Z���d�6�S�	��������s�M�˃VPk�C�;ZP���������=�L1M�����e<�*��09\��N��%|����Q�u���:��k�Z2C,cܼZ��3DT���{r��=�U��^6���VoՓU�'�I
��:����?{I1��f���3���eH���L�v�r��ly2`
�A�%�d_rM�O�[��4���0�+v��Ȩ�v�QI������2[�=���V��b���-�g��z^�I�,�G�Gq�{upY@"�����`�H�G�~�v�-G�W�Pa�}e0�hɛJ/1?�_�EMHsu,�l(R'C> ������w�#����̢��J;u�AD8�i�{�ð�?}��P(�@���K��UJ��e����~�Cr�s����=����8���}J���e���퀁��c����_.�S�H���x����e,�x�8�ص4�?���Y�3�k�.dc��m~B�T��f��^K���]�2�����qXB��$]��8��B±�(s�:%5�N|�C���2��B�[�{��;��&xn����m�B�#���&�]�5���QQ{2�*+1�n����lUp'�4�^�9�c9ONa≕@��	�T��%$�s@�@��	f�EQm㰛Aq�!��b6:r�!����MȍH���vǭ��#I�V�v��zi�	�sϑ�,|��8�s�O�	<(:�M����P�lO��Mp*�d�%�L���Q�c�#�!���;�:�å�^���;�}���7"%�V��z�C}����ɔC�^2�� y2u8�Y��"1\�צ0~����Ʌ�`J�Lm� �:�T���*��M�v�Ƴ������&�ey,k�R�5�RO~/�7K�L72�>�����LWW����i���N���<@`cVφY4d��iH���H�܍������+�'��qs��}�A��SޥNU�Qh��i92�J�^�&�S"-������=n]Q��E=���dҹ����$�g9���K#�vyv\��b{ ��Eyȧ������^a*zЬ��ܱ�'(����Ő��7~�1�M�u#�Z���P|�\7�Kjg-.��rR,:]��9�qCWRs���u�l'C^��T( �����'9���P�1a����o)tj�~R#��U��r�{X8�a07�������S��&��$���su�E�j�i�W��yW9��yQ�����5M@��W��m��uR�`�ʂc绛H,�ZO��b�d����2���Uw~��O���-)s��#�`�+���{w��1gO��T�e���B|4�)��Ӛqnti٥K��z;�����h��!���0�r�N���-w�d����
@�|1g����\���[�̆���(�L��W�-�� ���HcmÐ�p��>p�3�������V�k.�S��*.(k�'Ür�K�n�}�,�n���1_B5Q�z5s�gl�Mu�'Z���+eg~�!��3����it�{&�hK�C�8u{���,{���񷃊�����SYw�ZF���L\�Ĺ�\�x\ ^dG\:�e2��x�]�Нa�7��m, u2ق�\Sx]D�y��[k������+V^	\^���&�F�FGlUN;r�g��1���<��+�@I��t^�b:�^��M���)�����Z��D`�n�P�5��o��"��>���Z/|Ϟ�D�d�����tl���fC]���qf�Mz@���}���g|w��$Ą ,'�it�����|��4�k��'���������^��M���`t)�~��q�`'y�Rh`�e��bb�x��K�k�|���3`���O�������"i=�m�aD��N�tWBn���^Ѥ'���~5U/~��R<qޏ!>8��ÝY�b!�~z?�M:^�KSQ��Ûʦ�P-��6U�F��#�w�уL��]s��<��?����
n���@�'=�t^�Ȅ�ׅ�a��0?1t����I�L^^Ȱw�����?�3�������;�FO�y�N_�k��3�u�
	-8Y_�T$m�ḽ߃6��	������LQll� �޿S��ܔ�	�G<�səy�&8��#�kƝN���Pm�(����t��H���gA�s*$U��w�"�EH��k��!>)�X��5Jɒ�.���/�-E���1���s�˕�� ���S��e�*�F��o��D:p�����@�ЦŁ�Ob�{�0ߩK!?xu ]B�<�����G:y>���;�
P0����09��`�i��a���+q�G|h$2��.���L$WG��۫�ow~���o;�.�<�62��ɔ�ո-��iS��;�Cmh�p�Vݒ�"n���e�����Ԕ��e�#�B��{�%�>,By\N����.�����"�S۰��R�b�����Q���K=!�_
C~�7afG�/O_����b:0d8��81�I0�4t��L���d{j��DO���&��3,�f�~����qzL�;�:w*���6,ұ�,&���X��.�8���&�?5�p/	��"��y�s��}���7_|!�܊X��sh�NR1���6=!��)�wG4F2關x����[��T@�x͘oc����a�a���(s���<�V\ �G'�9Ȅ��6$η����	A0e�"%9j��h������_I�2���կ���<`��TA�B��� �v��ژ�w��v��Q�rO�D*�d<�
8��v4�g�͆I�r�ٝ�~�^�T�)S����n��֍rTKg�D�5�E�o�2�.Ǆ'M~(�>,�򓔾"��8d69�_�� H��l�f!h�� ��#�4Rp���S8�`�ڵ� �#dm�$�6�gw5$,���) �,�s�(5������i��u���������px�E[V��)����=b�+\`̋O�djN� �	6Y���߅�<�p�)5t����5�� D��!e����0�`�V�a,Kn���@���D�^�yx�;�u�^���~��xrx�Y�/��]fـ�Pm#���T����/�g��jJC���)jY���?o��RG��:���{��ֆ.<�u�)f2ԵZ<`���UL�sG_5XI7���
 ��O������Z�����Xp��7�Z�f����؉����&�ãy��tb8KXk�UtcHδb�y��+�2,�]v���,	�6���S�FR�E_��9z�i:v0���ꠊ9_wb�33��V
�IШQ?	x�6�3�.0b@#��(�ܰWi`C�<��:�._t���r�QG��_�¨O��ѹ~���L"��G-�mT��k�'olhn�;�P�_A�ܥB׳-긐�C]��cQ	r>&�7��Y���I-���gY�Ż�;UԊ�G f^�]���(�pzgh7/��� %��MkɗJ@$�+M�s`�3�؞��Й��(���BNr��T{��	^ץ��1uM��)*'��i���y����V�9��&J�W��fnݵ<nj��0C���ʇw���ѿ�NԔE�!�iT��~���ev;���=���/�eV�����Z�30nv���y1�Uoz7D>�5��������rC"����ω����(�lZ��L>��i_�_���ѯ�.͙)?��e�gQXw6�3[��"S�7�+�����:s.���4u�e�L��9
�x��T�������+k��W��Kf[��^�xp�K��К��`�Geqh�݋䥲��ْ�WaKE�j���B���j.c�
��*CM:)ו�X�&�e���>5��K%�EZ�ΐ��k��s
�\�_�^5=�(_)S�xsé��q���t�Y
��h|l��W�X�)].����C�p4��Z��H�&�z��^�3���c�Бx�E������=F��jf��"�� ���~9��?�, =��݁�0��@��hVQB�^�Z_4�;���O��k�X$�&��5�$��wt�Cg�w&��N1�+6M['%��X�2�pK�M.��8����p�
���˹ ��m��T�XOr��"�S�d��T 4Z��&���hF-Q)!r���a�<�K�1�W7v#�	c��v��q�k��f�i��XL����c��p��X�ZMn�x?�#;&k�2F[�K[T�.5��j�����8�z�&}cV��{uµ��/$B�_��5{n�J0mdFr6�
������ݐ�2��;�Y���J�Dĝ�C'퍖G�>r�+�V�)n���E�}�Wys�u�������4h\�"�r}�,*���l��k��N���vI� !033`�?�����`1���H�߸���,� h6K���>nQ�����2"��T�لBl?%+��b
���AvJ-h���>yH��Rn�:47^�4��ho Ԫ!>�ȝ�A)��#+�o���w׊��Vړ��:R�N0f^�ա2 ��X���{����@�ˬMe�R�7BBݝ�:�*��L�+������U�F��D$[�����"9�V2� ��zͭ�V��h�K��G_�oz��g��˱Ҍ"p9��րn4��o(�L?�lQ��",tM��yA[iD���{���l�h��o�[jz���&¦��ӧ���;V�?���Y7���x���;���A���2�o'ό��B"f���p�$M�%�vcX�O�4��o����&{�WZrdh5��[��y
���q	��|e +�<<7�'���p\��л�c��| E�GfK��y?��^.�#���q1
)�:�������CW�����ۓ��\(��!�
��5�5��Mi�K�[���h�������^��͕���A���4˒��0Xv�O(5I.����)�<%x��?�s��	��s�q���If�@�lf�T���Z5�V����'��[D�h�z��-Pxu���0�π���;F<b����aK/���co��z�)���#�T��L�՝.��a�
�^`��xPݱg@��L�S�����@�	#��^w�c�uyԇ1�d��xȜ��I՜��d�uKT�G$�>�Vf��x^~��3�D}���1B�֌3�OGK<0�Q�;^g�����|��P�	���=�Ôg��xA��-P�$�t7Sq��4*j�3��܃@;��G�W=�2+�m�������(+�4�3)�>��,鱶�G�'�%���
5��;l�@gG�3��d�jN5��W�h�ف���d�"F����C��_�r��_'I���Xz�u�9�F��E����,���`GmF���ˤ-���f@65F���g�|�##v�W����|\E���;��(ۍ����Kj�F؇���p����'(1�H		f�/�f�/����)	�V�C��3D<]Z
ikЏ����y�]�D3.6b��E��G��죙UΚ �#��JS�<b�I��b�ޞ�DJb���Co�ۃMpŉ���`�G>i[Sv��]p�y&�w,��q���k���~�<�#�|FA!���8E.��˝C�׳jX��{�g�d����,!�/�-�1�\�lU�0q�	�H�HaS�&㢞Α�U�"]���qӸfy��r8���c�\�#;�}"CB������5C�%�%)�B��Ħ�1���d<�@E�ԑ�٬L����S)�e�[E��"�o�����d��IQ�GM6~;�2f/�>'+yWH#�4��M�A#8�{���Ae�'���ؕ�8T�����_��$cȇ�A�ڞ�`����BT�P�f$7��P�H<�X���'d$��4-B��:ds7��M�ަ#��bx�����z�y}r�>��ݣ@_p�k[.�}�gҊ���.�dr��3N��]X@ �0o�������4l܄��PSDWѰ�v����uu�pzD٤D�ȁ��	2�����4"{�Ct��b>J���P�4 +Oʮ�%|B7��c*X�HT�~�'�� #UP���V*A�
�qA�� Nx�o�{ѐ��jV�b��t�^9Z~"�R>�iVe7��7�*E����H�">$Yݴ{�$d7i\R�s)�*`r���$e��@��L�^�Qt*�ד�uu���qa�*�	]
�[:���VcC�8kJ�zjcb�o
f$.��ޙi�� �,����ʉ���$�L�x��A���Ru*g�1;�7۵kR�Iq���L�wuOtS�ʽ)�#}t����!��9~��H�
�`)x����wD�6�ƌSRJ��R.u&���c�	�EZ7tҥ��ӄ=���h�5k��r�2���u�-�wc}��ä��t(���\c��˘�q]=�B��~Xc�	KIHĬ����:ͦ�ib��2�%�-�l~�>x���d�.%���.J�V�ؑ�V�S2G�/����$�ʖ��H
�3��m���f��t)���F����Ս�a�zu�'0X0!.K%@].50��p��uat	� X`�*�.�����f����_��8���R9[8W�89үc������~��C��M�_�Ɖ��E��,ew�O�5��"���Ε^V�1�K�XWG��|���'��9����	����\N�>!�+n�4s��Qa�I�=��k�4U
��d�ץ���)�bHA��ǣdNZs?P8���a��WK�c��
�ʱe���:Q1�r�����^�24�����"�XPꪈ~��A��XG��_2Cj;H�������st@� �VkN�20n�[�;Hd��dsuK�ݥ>�R�Q"3[	ן3:ޜ�U	H���q�#|L�Z9�PVmF�߬�0|�NH��]���.��i�(�6+䍤�d܁�A�C ���+9#���+�&�@�<�thZ�>M���������[t�����'�k���S3�a ��K͇jWRW��r��o�/Tx ���q�vb�0&�[c�z]�������y$S�lC#�>腞�4ޅH`�����0�覄��'^�\u4I�C�g�wX�lR�j',�f��*;>UR#w�ѯ�Y��cr躣^3��+r`!o�Ψu3˘�(&�rj���v�kX))Jj���|ٿ�l�gb���s��elO�g����c	�r����ٱ�^�w�΀g�캓]9J��U�!�$y��,���NG�}҂� U˂��g¬�۹ENП�'� �8�|�Ъ<Jx�wӫS�~ݯ>�=P�1�`�Đ���Z톧d����/;٪m��plr(kn5U:�E�N셪��lH'$Jٜ����d�Ns8a=TD�`��^ k1bY\	ش���.��jp����"ۘ('E^�	�+���\03�K�Ã�HM�U�Uv�8�c���!/ee~��%8�
[�����Ti���e�%�wX@1H�ۘ?�eY�9U�� ?���]7N������l�0F�x2f9�pi���A���W� �����m�`:!���G�ȩn��F(���i��
ɑҠGBw�����	�{A$J���H�>-�"�u"��z�ش��D0�j�)��keNNj�5���B�b���.it߽#�<t��;H�++�	�p�L�A����6an(�ׅf�p¢D��}h���kop E9��z�;R�P$��V��
'G6�����Ӧ�������y8���y�TZ����;��SǮ����VQ��R�� S��ä�y8�����@��y\�:I�~0v�΂���� �'�:b{/[�Q&]	;��B��$O�H��ej��	P#��@�+(���������,��+�)#��MQ�?0 �N$�"2�B��ƫ�T�+��w� RQǷ�k!�����࿧@�(�g��>c��n����������%o}A�~-�] ��QZ��P�`[r�j�h�_��c�PO$��p�_�\."Ĭ�BcS@�م�4�?���/�� jGD12��V���Kc�%�x�D#i���� r�mT�Ϸ�Kl%M(NFe���q����K��-`,&8���1/��6��(�[�]Q���٤{�xa\6��XB7�6Zo���u�|���G�a-����|�BJ
h�����,�m�������{�Ҷc���qY�ͻ�4� �c�gS ���fXBp>J��ak��{�l�0=cL(���V���E�g�!*���S72�-X½��S�J���.N����M�I�螈f��-*R=h����*:�O�P�l՞1�=/�4E����qUY)�9}O2����$�;��~�o0�SU�:�r����"��aB��%v�ӈp߰��(A�a��XW`��j��ݫ̣�u�}��G�[��8N8tU[{	���}�i�/G�Hk�tR�v��&����Y{��	���Þ�6�4*��aU�P�k��|�X���q�>c�44��N�3&�H��B��v64��Kc2F�t<�a �d��e��Mv�ZE����c�������z���,��$�bK��(e��e_���(�+6��R�:p�t�I56�e���>I��J޷5o��:��.G�[n�1����Ɔ"�]tk}m��V�^����N���^��	�a��I_����6�����;ѵ�6����a�}@ �RDw?��(�G�|;��wX;.B�]�*?пz�|H�����m�ߺ��E��T+=�X&e��b?mD�3��E@���� ���Ծa�Ϳ��n���y�G��3cL��1o��q��5 ��[Gϼ_"ܾ���̩Vx��.}7FAJ��pK��td���u�/ʣ�ޝ�p�sN� ՃD��S5W!�/��:��ޒ��s�U���ݛ��O�X�%P@u�F���ۂ�E�P�@fIGq$�O����Gv�V�q���XY��D��a�����,�k���<���H,�w�5��U�-�8lA���U��8+${`�[���K*Y�w���hd�t�4��v��S��﯉0Ykw2�NT�4����!�*?eɺ��1�N�?	"�'��b�;������G���'���z&Cs������+/kݹ+����m�i���񨮃��c��3�|?]})���X��&vR��-�8D\;œc2��/&Sb��꥙�2�=8�r��~���4 bqt�	Ҝ��(��� C�_d�	��(T�j��I����GKv��)�^�y�h������P�#��Բn7/����q��~�����l+����rqU�?ən��Gqߍ^�����9��t���Y(�b����%���6b�Sˑ��pSṼ��Q���Nfڌ��K�i|u�״*� Hi��~?��Fo�+ٳ�}JC�K�����,�tcŁE��죀JͧXR
�B�	���"��s)-O�v�A�Ĥd�g� ��EwכC���ÛrV �lz�b�>�er���|_�_<�r�����1�Q�.pĒ$ہ���,}�:�1$�QJ�t&Wh��@��~z���;?���\ PIa��/�evI%`�ԛʝ(Zq#���
��bD�޶(
��@��)6�_��7��X�i8)�(�T���i3,�x�F�D�n^�����-�l��Xz��o-�D��c��_�Z~��Z�v��|"�B�����4�y�ţ�D��bͮz�팠W�#L��,�d�n��у#������.���ӡ5ݩm�� ygG ��ս�����#YX��X�c֖*wO�#�����2哃��\��)XM�pgjIu��|P���B���@M���
����-��wJ:@Y��m-(�u�����#`�����ր_z�ubs"�c�C_���Aɕ�;T����$�	�C�O�`��`�:S<W�r�j�w�j�z8���8ð��'Xa���h�S�gy��z�L��0dA��dx��VU ۵�l��yq����ע1���n�u�HNP�JRI��|7&�,S�,O[�xF^S	��1�)MX��/���ij��i�u�~��Y� 	w�1�^�|w��8T˪X�?�RA5o��%�c��W��i�t�A՘^�GǬv�xm
TC>L86e�{�n��P}��^��FCh�3�-30��F�lz�� -|e-��N��d Uy���>�
5��j�∮/z�I�Gi�<�Nǧ�����/�es�i�*�!;C�3<|�DW}^pr}`�'��8�r�Dnɪb<j���hi�|k��ȕQ��S���b���Ȇ`B�AW��ǐ �,��/[���Q@�p��D"]�G�x�Vt'��x��2ok�0�2��'���"�ÚXg�N��&]��נDs���>톳	T��/���s�?�;�<_w��gŭOw�-��^��#����-�_D�1�o�=�y ��%':��>����'��9B�V˜�;�&I�k�w���xs��"��v{Y�Ҹ�V���𐬱���+[����Q�  �cަ��䰍w�ͼ��ڔa�G�[�Rz��菰�7,���]t��.��愥ן��F��X��_�����B��>>��,Q�[!)�7I.(\r~PX����8�pX���M�3��Y�����5���E�jQb�ȟ��z�_��\��R"�ER�������˭�+u.{���v�_U�5v�2�7w�Mk��!��6OST�[.b�}�,���l�́śu��=[�^`��rg�4�q�?!�
�Zadv�k�@q�9�3��!.����V��1���H|�(�+�#5�ç�{�q�pٟs�+��a�O�]��^���%��Q�ͧ����1EU�zM���tZ�\DBDd7�sC�{��S�cm� ��0_ �dW@dݻ�坺����b����M��P$��<y���^�U,�R��Jk9���׍�nY�3����żTg�M�iSPc��V�h���Ϻ-�u�P�)�aZ�7� �3��N�����N�u!�n���!2���g=�S�p�	�T�8�ﭕ4f�=���>�\�F��Mz?�U�Zv�V��$&x�<�N���6k(Whz�������}B�8�?hbzT0A&]��!�aw�O��X'���N�C���u]wb�z���w+�p�Fj$�q7���ț0s�<� �{�ll{ɟ� �gJ$���\'yظ�J�'�Mx�w�����k"%���������CA{�
�ŋ�iG}�*6�Q�$pzC�'l�܄��ワH+5�o�Rݣ'Sbo þ[N��a�Q%�멑��-����Yw�D�����!����2vn���`�w��j口r={��iZo���Ku���soeĪ&�e�|� ���'TL�R`7f����Z-����b����(�3�]s��}|�U��
A��4�u�����gmE#5Jc�b��_"�!��c������é�Q��L'�S�@ǦFƺ�-ú�]^��]K�g)D��sKJ�. ���	g]zX�mV��@��hUN�}'cr�TZ0���a�D�PK�h���x��i���Tf���D�}R2:̺K�$�D�X#�e�����w�=�����v� ɨ�ζT�$#.U ��l�������,+;���1��.O����������qx�:���>�;t_��ȝ��̓�W�`�# �I�B-�Lu�	��JY����6�T�6M�[pr����^����K4��.=۩O �0ޏ?���uCC��
{s/GB�LǄ�k{}d�_%�P��l�ڒ�:=��/���s8ғ���1�i�3v���W�^��"z		qI���r��E�)u��'��sz`����%����!���TB��>����b��� �sD�BS�cjux�&��	�0P��"v
A��g*٫�d�����}D�<��8�_�Q5�t!ǵy�q9���#m#���M����X
xË��)@(,}"�Cj�~���M�)s�� �GH�.��e��c�9�����`��A&�V48H6���V88
�Y���>6���N�����>���9�\|�]�L���j@����-�\߃� ���[�)�A�����yx}}��Q+�d;H����O!{h�4>�L%�6�$�mn����p�q�d�u8u�\&^r]�ҥ���p�"���x;F�\�uv�㮈f ��^h�ؠ�˥�uM"N���W�GD����ד��[^��H�|�#��bp��S�����(We&�j;f�P@tɒL�˼X�.�����ˎs:~=;���ɒ��S���w��_j�e���/W|�J�Jc���@��y���P��5
3~�}����I����~\��LT���f��F

�ğ�&$���� +V1vo���T9���?J>5� "����]���Ā���CZ�;�v'���Hڅ7�s�CvH��ߚ�֤'D�AHF\\�W�8�=a����G����nKZ3 �#?��yK��3P��Z��2K�HofBg[P��[��n �N���.du0�Q�c�u��	f�I��c\	F|�op�F�o&h-�2&q9�����g}g=��;�u�TC�$q��T�ez78f��DGL����v������;�e�!�P-�D���V<���l�kKz�YW�&�3JE�������}-��d`�!2��R~����*�ѩ��(�� td=MR�R�����l,��.0"{�ж�f�Q�����c�fc.a�0h-�`in1J&P�E@1dw&�	T��x(:�u��Sr��s-��D_���x#3���Ce�b��!Y�x,���k���a��"b�����g���v�_��"����;�Oj���W����x�.d�$�����;�-M:���J�TEe��<�\䳄Z�����^��ܦ:��e8��0��-;X��ϓ��DSXo[6� 
�JP`�|+x5�S�vؔ8e���� ���h���;��՝�s �:վXX��j�Ѱ���̮�$; ļ�n�΍�!\��&��񜍚�$N0��E�K8�d���ۊλ����xm�-�v50sP��t.�&���w�i��B�s��KQ�h~s���}; �K��
��mR��A}��Fc"Z���"8�nL0Ե%���=Mw��t�Y<{��+��V��%3�o�e�wS
�&-	�@=���ᅧ��j���� ���T0]M{s�I�Xa�K���V0y�#��2xq$������W�cwy��*���c cq�?�h�|��@O�������['��e��A9���x&������� �%{E0�z���\_x̆�]���+^IEp��;oj;�9���X�<������X��ϖ�8�z�<��M`=pn3�&rf诋��e)U�{�!��?A0�X�I�im�&�Y�ސjZׯ��)u�¾�y�����m�I��uᄒ�6X2�}�H+�L3��|�8�?S��7od��?�Vt�{��7ݍ��u��Ц������D��bg�V�XbA�^ٙ6i-�9~W�P\�<����mTF..2�E=�#��ġ/`&>OO���,̈́P6ƫ�`/�-ep1��>擶�Gm���� ���ȐJ��y���G#�V]�dRӂ��:�4RT�6B��F���+3m��һ)Hl��&�Y�괷hY�x�R�7jA��Y�{�a�!(�l��v�UL�������kK�^6kg�R��@�N����)���՘����R2��gCX��I�B� �	.3�NV�s7�έ�C��&�΍W'ӷ�f�PFS��H�����{Q(@���>:k?|���������Y����K���S����ŧ��A�O����5z�1p'�|�bB�&�J�R���sޑ�@2Q�X�qAN254��-yL�;M��{T�f����>w~Ү�^����;��~��!պ�g�/�u��"��W�G(b��8p��Ai����^=8����~�r�#	�ɴ�D[n|\V���yE��:A�T����i�2�:�Sd��1{έ�9�����%��ЬdB=Hg����9�b�w���P�AɊ4�NC�t[�:��t7�c��gfcx��ub��v8E^��_�%�\L��AqD$��*�\#�@#��c�S�$8�3���5��,0�Pʾ�z�5n�N�gGFc��N��)��>�\mD����#��N����E:z�@˽�RF1���.l���kK�ʊ�5��ꯇ9ʢ�<�_�C,��c�n�)�a����2��_�ۍ��ϾdX*�jv�o�m�`:���	?��y��3$K�։7D�v�|�nT
�L��m���2��G��_`��as�|^E���èu���nAd��]�<L?��*��K�y�b��N�C�ᡕ�F�����]�Y	"�6$��<8��$��z®J��j^�٫B���8�
h�XSN���x�R�&!�}�ѷj�e��AH ԡ�@��J6=��S<	zK�`{V��R`���Z9�N,�ދ�q��uk"#��@���F���X�b����t��Kan�G!{a���0pTaIRW+�ն&&/�(
���`�l%c��p�-1!���c���݄��=�q�U3��RQ�a|�&_&����	�j��1��l7*D������]WW�Vj�4����������,=��f�'c!�+���1"�1!��<E�d�z��;/�
2:�R#�,P�\�@X�D��b�i6����S�\�r&	�6	�dk�F�j�|��@7',%��^[@TӇ�$�8T��Iɿ�T ������ކP�
�s�k)��	�T�s���1z3#c��U��ꑣ~Ȼ�:����Y�1�d������_"�������;a�q��H<�w_Y�Xn���A�v�Zy���pψy^�1vh���7�&�E_���=ce�Yi\Kf\S���������.��v/��MW��샹w���D�C(�p
s���)j��mB��n+���N�x�;J�>�qZmsu+��~*�T�Dt�B������J���3+Lb�O ǌ��x鄂��ԅ{���竿�����T�#���&1/���L���� �<h��<qpˤ��oԼ!�S*�m�`M�ϕ�M��|�4޲�{Z]�~�������c��+r�0>h��\C��癠��li��Q�$��8�]�(��S�nܿ)�ɧ5]�G
��J̣��;aԹ��7f�)���[��B�{��0>:^��[V���=f]SӪ��.�����v�E�����WP�_ۦ� �O�E��>�*���:N��옹vn��#Q��}w�%�l����Ybz��4c��t��b8��lOJ2bj���q��Wx�T�����Nۺٙd:����a<�	|p����k�H��Ti#r�d�O�pd_�g��c�Xc��iS� ��������<@L��w �_��,K�[�`�3ޅ��~k�#�%�
����\��De�����n�cE�Ŀ,6�7��� >��0��t��Jx�NrQAf����SA��j�z�-����^0r2π��������<l[��0H�ǿ@�e��Q�W��_�9�WC6��|ߝSp�W�4�0�i]NU�>�j��.�Q!S:,|�Ƣ�c��(\k���Н��g��B��*�ꌊ���[�'�����߼	9 D�V��J��҃���`(سC'�A��Y������Q�Z��g"Q+���c6�0�-ހ��U=\��l�hno ף䣇��"�+����E�ZZd91��lH-�k+�m��)~���9��^d�S,s�䆜̄+�uꑤ�l�~0�ؓW`��b�N�W��!,�#F�7�JEu#��_�)�q����s���׾�_a{FA;yh��(����0�xF$! "�A��'K�y%���m��}�b��kOi�+�%V;4{��~e 8��%\�������5�e��R����b�O����tr?z�������g�[608z)�#�S���/h�W��?�{�Ňe-5��ҠJ�� P'V�z���M�|����̕�f]�!Im����!�5E3�Y���ΥԠ�?E�M�4x���,"�����l6k����p�K�����n���o�<�� �e�p�� g��Dt{3X֬��u?�Z�n���p����ܣ�q��{B�2�T�+Q�]�qCRȠ�>w�����8McY��7�,-+��,Z�d���\.I���n����!�l����2>��F�"?�->&���q:.����B���.z��HE�ʗu����5��F-���}����$ln���
�]�Xs�q'D�7�@�1��-��Y>d�Ѯ},[���}��������8���Wm��z��A
P�ݛ�W8MA0d"��H�Nv�ߩ|WTh���[ZR�3ڏY<ì@�x��7z�AD�H�mS8�SOu`���4)��6PT��f��9��Ǧ* #�{�Ҡ��<�;�l%苛O{���&�����򹵬����0/�����C������Q��C�_�DP������~,o��o�[�]�m�J�z ��vT\��O��U��+,��G׃U�_����0tW�U%^��Fx]�N0�����Oc!J(/�L�pt`��,���nZ�!#��qjm����1I�1C�Du`p����s���E��3+��W
U�CO�,���щ/��۝_g�����l�<o�����fӋ� �A4�..pŎ�)k&���H�l&�kH�$a$���r���rpd�����tʭ�A��Ɩk�*,l�h�ǚq?����3�x��L[�������c#���CZȩS�"�^��'�ܲCɣZ��}����k�CQ9Y��4�<�qQ'u�N�\˸��d��Ȝ�\��n�w��ן#�xTl�,��r:���9�%��9��Ԟ����2�"8l?�A� ���U�G�����ct�۫!���\���(u�h��2�5��Z׮@�r��Ų\�A�f|�~�"bm.���K�q7�ns�6��?�K��.x�p8�s��z�(���13�$x;E+w<�N�L���戨*JUY��"8w<����@%�br��쓍�$��k����P�Y6w��4�%xB�U�k�e� ��O5�MO�Mu��-@p�f�wz�^�@�ʨb���a�a���� �	2���8C�rN�+Nc���)��������0Ev�w�Wr<&-���>��+����;z��JR�A�d�H��@��Iq�6xo����qg��ȼ؍C)�z��h^}B(nL�����b_!H\!P��5�W�Gv����	@� �u���J��M�t$�d۽s1��t�\$[ບ��Ӳ�ǽFRq���y���t
^�\+��f�č��V�!la�<t0g-�� Zu�֐�=fbv��ꯜ�|y|ڐI�zƤ�*PKS0����ԻȘR����Rb�w��~��*EL^�Hq�5��ὡט7⻳�'�k�L3%r܃������$b����\����?85L�ދ�m��<4�n"�S�!�����n����oƘUg�`%�A\U���(Z��~��i~.Ud�b���[�J�)�H��kړo�
�6'#��&�e���'�ǂ9d�H��14+����@o$�֩�Q2FB� ��h{����%0��1L��3�
!��2�«�9PCM.~:ɔV��6�����*�:x�E (i�\�N?��E��0y�j-[E�W*"���%ψ��D�m�>�K��SR$��IY�Bj�c=-!����6���W(�����<��9���|u�7�s�҅P����%�J���T`)��|(а'���2m�~�b��"�_W��s�yM�3�����X���On~�J�6�F���'�X�R�����$ϧ!#cU�$�N&�rs���+F���)�Ԡ�^�ʭq'��l�o�������Kj�K�%�̕m=�<���d)�� ���r��BZ���=�y��pU)���ѕ]2�N�z��A1����~�m�n�ܢ���7&�L�6KU���GvJ%���^����$hh�Rm3��\d�:�Bѫ;n��H��.ݕ����wV	9)aDI�0���	7Bʿ�/U�F|LX�5]��VQ�>�J��.j
������j�!L�Ed5��mZ����q�/��d�V�ӯ!4�(��^�S4������O���@�8-�*C>��|�Zд����ٙBI��k�MNqΏǱ�;�(BM�O�?o�|�1�~�����u��c��\�[���@$�%��v�r�p�&\�@�Q��f_0���z8���:�z�9U�%�@�To��aL!"�F)�������Ђ]���EV�L�u �C�;��.�7J�+eC+n���L6杒�WA�T�Y;įѸ�9�:W�������<DpW�g@�S���As��eR�P3�~��,G{GZλM��Ɓ�A#Ƭ�F�`E.���_����~~C��4[�W�
�����&NR(��EBZG��3@S���(4e�w�cA�}�2!���<�Nʘ�츌>I`��s"l����޲RL����HU�����%��*�î�I��*}� ���Ae�t�S1��݁���p kt���� fb�6f���S�9��K�(���@����+�`X����R'M��!�����\H=�ͷ7F��}0>�. ������Gr}ް��p� v��u�E6��l\��'���1����z��$/��Ե�gb./3Y�9O�~���,����"�;j%.�ԫ�G��aƐCJسx*J^Q.+X�a"�>��8�U��/s/@q��~����h�R�*�æ��M&"p���$��o��	gϯ'5m�->��=�?0���b���J��1m������
�dK�����b�K"˲�����m�[-q���#���yB��C&�7l,,��foe�V[-x���[�	t��Ƚ}�|E��n-�6���qB���������q\�.ÞZ���Gl���O.G�ug(���w�yBeB9��?��tГY�.�N��uhy4�~=A��	a,��P�}G@ �\ �*B(z���Er�T������(א�N�FP%�K����nrd�\��u�>�ٙ,-E��y�R�������PQ;��v����N��2/�3��`��([+�^aܗ?��|�;R㘯~#��I��jb�uCs�+s���S#�՜���ɡ%�-%ޑ�����T���j��(�ZApJ���7�zrS���*�EߐSH�_�FK��g�j.Ξ瘼�39���}O�Y<�4���T`�d���fn';�/O��ݩ��_\!J�����k�r[t�����U�\����ٍ�dI&8����Q����N���4�'=�d�	�dp�I���_)��+\nqZ��׃GH��7[
1��K�Q$d�oA�Fe
�@^�Q\ߙ�u�F�=E�a�<�%j�)���A��%I�<��J"���7&|��.L$�����X�s#��ߜ�8K$Dr��@n	n�;�
m�nK�"��?�6XP(@��_�P�'��m�*����g=jR�͝����
/��'�Yjdl�h4�cٯ�78,#ё��S��ۙ�غC�,x\�H�����C6U6�.�Q�J1�ֻ���|���YP�V����k03Q��Յ�>�e.Xwo�Q2��m�J)�kU�[z��D� P��-�utVc@QG�t ���b&�9��_E���v�N��$����v2a�.:�Z��!2��"�٭n�J�cc&�Xv=����ʤ0B��;6p��Z��:�,  :%c]v2��a�W-����h�S�9�X�Y��jYb�C[���t�s����S�0(���k���,����x�©`�Qk�KPH��2�ȟ��6��]��)2M��yS�I�jfNpZ�ry}ӆK�/�r�2RBm�˴A� C��c�W��E���`��H� (
Ԋ�V�hJ;:f�/�.`�t9�DvY�?׮l+{�[dg�vm������}��aw���ZPy�����E��DZs���{8�:׸��Ђ�A1�ͬ��7mM�� ���
6��+ ���D2 8�o�!c���r�G�`:�}A�m�ѳg�{�M�������F���~��cM��c�$��f��0���RG����#V�!B8�$&Ɩ�v�nE��I���Ɉ��;�}`�����p9M��E{�������T�~���y�]��f s3[�FZz&-�Sͭ�$²�z�Q������K���\�?��Uq�u1�`�d�`�S���	��Y��{�3�v�5/ �.�����h�.t� J8r���*��H�~��ST�..۪��!����S�����T��Q�.��M�E��	9oR�l�zj;M�띂��:G�K�ą��0,,�5�H���;�T��4Ï��vq��~��<>��JE�Ϝ�h>.�hK����/YW��"+ɗXS^Z�i�������a#�Nc����xUQTY �p�_ۤ�Sz0��h�.I!�ޤK�T2{h�o���k
�Km>X��S׃�H�v8�0R�.�5#��A�B�G5�������ǋ=g����^o�<q��@j��8�X�tE^����L	�:�<� YBw���
��!��ju��<�ԉ�Cjp�}w��nW�W����IQ�mSh����{b
M��H�(*��{B�V`�����(�7�Y�D~�hw�e5����8ٖT�*6����$5�h��hV�i�{�^��|���8�T_)c 0�{1���/Co=���Ԭh���ޛp��ঐ⌲+��M���4Vi�F+��֕ҽ*6!�)>w����Lz�0*	!��[�w6�\��(�=	�V(D�;~Tel��o���U�?��gȢ&s�Z��r#���8Ax����8�m��!KO̩��O��횑�����VS[��Da.'g��tM��C���K&�����W�lIB����e��_����t�
%����J�*��2 3�?BF�/[�w�2|�n^��1}�N��e+:��Mʤ``B�e���a���㷤cM�f�
)�!7]T�O�)�ō���Zj,j7}ߞ��}�xc�4����ag��I�Y��%�7Z�W�� ���� �9�e;��d(a ����]A�m�Y�〤9���]}���§~�])g��0��%#$����8y� ���o��?X��j>�<#\�'υ������M��ws@�n��!w˅��E��S�4��8y���ÔS�*x���R���  � <���!ú�B$߱Ā���k�[�j�s	 윅�#��х?����z�n��tI�B<�tV �5uKvL�.��*�
��;;ᓫf��{�յ($Qs�e�e7#`���9�Bq����� 4�7"���\�� ���e�]=� �!��2z���V�aU�����]k�R����轈Uu6�E���l;9� C�p��X� �.̪{��?�2�!a�>�nyr@���틵b�f���[��T؞,[��gN�ҠK+*)S� `�y����'��\��;}���c�Sa��P㘆�08��P�����1����ݎ�l���c�<u�����w������}�XڔT�?�X����t���O�پ�_�9{]FG6�����X��>bw�n/PNZ���>eA�*`��s�����r���w����N���0���S-vdQ	>��{���x0�*�9�3��>�(��j	�r���]���͑��֜K����f����ZvE�bӹ/ʾsa�S�L���+�<J���a�ec�����p�f0���
!�CdH����!SP`�ԋ9��@HU���s�B�gq��~޵�޲�.�"��ȼRBW�6Q��npԸ�$?�GmT���W�N�o��y{������(�G]6�J�����S�&�xxP�u�HB�и!P{s��
��mL��d���e�?o��u`�cc%7u����j��S�`�
�ɤ�I�(� i�Xb��F���ŷ�$��xfo��:����쐝@�6G���:1]6c�<�ۑ�#U`�8�i�Lq�(`n?�:�_(U%L^������7g���կ�~�m\��l.��ϴ4Y؝h��u�Q7q�Zh���X�����r�(P���dh�Dh��t?C��$�E�PS�b��m�
�$���Rfp%��$NM���|�i=9'&%lL��S���i^����f����L*�h��;�ﮥ�A��������;?xG4g-�����G���+y@�S�����~�LѾ �x␧�I+�%>�W{��قt6K��Fr]�������=	E}ϩ`:�Ԧ4�I�*�uκ����'zk��-����X7�}�\ƶO{El�DK��{.8Y2a�=z���kԦ_�[H/G�Sbb���ra;�+�A��ДA��L� ^y~�Nd�4q*��?+�&�w�aH�-�-��^c2유4�q�[�&�֡r3Vw�D5OL�*J�f� �ӡ��C��n��b���0��Qm�*��E~�vT�]P������ (bN����Ow����z4�!��2c-��P�ƥY~��` TPqUGsΡ�����ɣ2=2�6�,|/N+�m�2۝��_V*�"P,	P�V����ۘ�q+3P;����E�	��%����v2te2C�S�_������_���/���J��Mg���նY�ۙ�F���%��7�'^#q?�,�#ʯ>\
:0�cvPzaX���.��L���"�/,}�a��!<��#��xER��|��Ǖ�
�p���˭Ҷ4��|۫�RyR~67Շ��\��	���T�"Bu��P�u�+'Hw�i��Q����U����h��R��j�d�M�T�Rc��/��Nk?uH���Q۲�g��U'4��O��&�?ͦ����3�p� m���J�4 �Gy��Të�`Rs�x���=�ݩ�CD�,�GGf�!�ޱ6���I��%�5<�QMلj���t5\�-\ '���))b��:)$&�>�)�"�M�m��I~��N�&y��T
��x�v�o���=�-���}���u��������z!#��yF]4�~NN�����+PO�AX�{�d>4:,���\�����߀s�io�՗4���-
,7�Nu5n}�0y,0*^��`ݛ�o��A�A��[ݩ��OT����S�2�r��������W����-�?�O�l,]�U�?@���V`a�F:!�
z�	��f7 �w�9%�y�A���@!n��P��ز����>G���ǵz�2��S\mtj}l�g/m�@�t����S~���%Ћy>��ً�cl�5N��Ik\ �Wg.��ç�A���U�L��#bN�w�V�d
�X�L�9v��7��Zj9�h���BZ���"�_���+p�;�$�-����M~s�j��,�����?j<�x�®F��鷧`�F��?��I��	e�x���O��D�~���o�i7���E5:J9An\ʼ($��8�/�X1�W��m����m��h�30��_�y��g8�N����3\jg*W&Y�"O$=�X�%��9��`h�J����2�}a��F@��sG�VC�H^?�'e7.!w�2[醬�u{}6�:Z�}ro^��/-�����6�yiݐ�����L��j��{�;�T���|�h?��z�Z��b�@��C��"�V�Y�>l����ܟ��\��*pNs�L+ӑdޫ:�Y-N}���B��M���m�����CB.��P=�u��<��l�1Mz�����h�S:'4RJQ-�j7��P�>�E�h9ٺ0A�ߛ���=LX@sO�2�cy�>��)Jo�����k3'�eM	�J,D5��qv�����
r3�ň^
m��y�����-��5�t�N��+J ���0�Q��܀�vs��N�+��s�!�J�weN�v��3λV��4���jV=7��/?�lH��oG @���G��2�`;�\�4�00�9~@������v��6�������\}�>Rh{���>�V͓��<aI��ǫ ��o�Ԗ�h�J��̷:��z ��s.�md��ze:� �M}H,lԉ{�O�60��Rd���1a��8t��и�&+��nO����ߵ;�X�%�U�iFLu@����RjM�KG���s�R����v�תe�7�-@���t�\�R�T����D�����gV%'''�K-HkFI\j4u��7��+��ŎR�E�ޚ��a����>���o�g�����|t~&�.���/�xQ��dJ�	Yo��y{��:q��v�9�����I���ڋ�kk�|G�f��� �i�9���t��e��n�y�#1��<�r�� ���?�;\��w�a-/4�)L.C�̒f�θ����󧅚���d�Dv.N�6���3ӌ3�'<ю\Ka�%T�j6̽��	�#G�c��]�( ��Yj��E�,���A�/�Y��z^�`4�X4 �K(M}��Y?j����4��2�'�`��D1�i���	�
�|�/>���uT1�dF3O�,���z�ZT�g��cib��d��2���P����f����b�qM�Ct���	�~�/���ҁ��*Ya�P��0�(!�@�-�\��~�Lu��$D�$3���5���qR�B��M�b�2��6�fjH�uJ��3_<�	��ΐ���sl���>�J��|C��{וB�q��dH�5#�����K�����̍d3�\M�q��ټS����ZRa���(�@�ʣ:�������{��aG,}���Y��O#���0�	9W�ũ&�InF���7��AWc%�f�f���e��cM�H��f+m;٨�?O��*d�d�Ә(�~jH�#�r�.����-�yÀ�ߞ����.��3�=1Q���;�S�m��R�g��R��yud	�gE-,�4Is��y���c�����{c����8�}���b�~��L�BE�]�XT�������1��-� �v��{lIgs�l�_�snk�}�����O����|{�E%A����;0�*փTTN��:H�aI�2�G��l�PҒ�ֻ�(!=�o-^�C@InXM�p�x5�`w��lL�1j}�>�E6U4=��o����4����gh%��K�PHhL��PH��^]�Vx���i7��Z��O�%M��M����2���WgI�!��K�Ͷ�{�>�C�A�� �\�gg�dn������*f�� T�����Uk�L�A�l��YAٻ��z͢%��%N���xH�� �`���>ہ|���F?M��Y�=��uZQ��i�%�D�mn,����5�߿[z�X��J� ��$�4m	������8�|�xJ&3�§�L��5o�����5
��`��l���C���d>߻��?H%��-MA��&��U��٪�_�q�B���5m�oJk�[lFz���ɦ�Me�=��R�9��I�%T̮}�]x�+��7XH,`�Ge�ҩC�Mmݠh�r�q�ff��V]C@jғ	�~�7��88WZ��s��x��=x���j#u �D@K����Ƕ��wG���y�c��Z��3��L�Q.�t`ҫ�p�ŏ&���rqv�_03�=��c���l�N�Aim�
a�������V�U$b��O�/�w"N��!FL�o�Yu�1TTj�F���/`@D9b#��*^�I��������&+\v�Tz�fg��zuNI�8j��̯�~!�5o�;,�Ci��U�-�R����%^�}'�/�+d9�f���3�B��4o��YcΊ�dH�*([B�[.���?^j:��>�dm�i!̤̘������!6����h��� QS3�U���3��;i&�0t����5��eL�Q園����#��6�iƫ�/���5(�͵C�1�)K&
U7��vE|�Ce�j����}�>����)T��fU�OE�)G��{�[V�@����,����G�8�̜��-���c��L��Θ���b@p5ey�1��7���pDf�cwڬ'�%�	�>d��Ep�*͗nDb�@D�J�K�:�$.!G�Kڙ�lRW�)zN6@����%G��&�*�n�fE���7~2[����2P ��M���#��r�	�/SIx� %��|[�m�t�j ��|y��I�,�vA�>Z���(ĸ}A�khG3�{dU�|Zb]4bfZ����Y\�|tk"��(mtǹ.wj#N��\"�������^-�"d�.6��.yN3i�)/!Yd[���'�#�w8��� *�X.��7��Vٻ�m�t+ul��(vm@m�7�+��h��7�W���F��8��z���:�V#|�}�X�ܑ���'T�z��O���'P2��x���C��� ���=ٷ�Z�����{&po��7�\��+�UR��\���rzq�>��qS��]�joP�%�p���0{��vMu�P�وC����=�l�7U��*C/q*�Yqoܮަ��x�rc1��Y|_nX����[��)�~s��̴;=S4?��^�6�"����|�h{)W\�=�ˬ�G$�^9
�tU����`ځ��&��(�A�|�R�s�-L�n�ީT��ŉR^V�0�`)D<��38q��1�Ѝ��M�!�؁/j����Y��pIP�F���H�@�g��KC#y�poLK�PEة޲+ ��.i}J�be<�#|o��\�8��Y��`l`o*�r�';E���l}��V�C1E�ѱ!`h�<�:��n��ac���3MU1���]l�z������O�*w�/%��Vo����-�TN2�+��t���ưҽ`s���q������$�;��m?+�n~���jX��M�¨yv�duV;K�����������2ي k[m�-2���ļ�!���Z��!������xl�)Y!��
Mh.JlM��$GZ�?�k>�u��C�h�����s���]M���� s��q�l'�Fm��39�'�P�|:V��Pz9y`�"��@g�h�뮼�K5Sa����ZIA��c�b+F�@�D!��(wlG��˧ǥ��K�Cz�Jt�GAH�|�����������>�s�w�@�p�6�!���11��kk�I�ƶ~�,~�N�
DG���;��L����?�M�����P]�,�[��ɟ�u��|��S�R�'��\uiR.��o%V�0e,k�C�C79�W�c�}��#c�˷а)�/�:����L�^��N\q|���V{BC<XS����PW������Q�4`%a2��w�y(�cA��8^)]Y��w1����_i+9�;W�)H��U��:�;���$1�����-�����כ���X�p�[�8�
��h��7-�kN^</d�� ��70�������8+R%�S�Jn/�G�|�Lw��}���J���)�W;��'���o�kLh��jز}C�(��Il��h���� ]��Р��17�������Tٚ�>��h5�"������ւP瘟yX�����uZtd0��_����h�f��s0��9w�*��}VGo����~�����g��&���7�1S9����4�Uu{	0���c\��؛�������+̆0�m-%?�l���{<ѯ��,/�o���2AĠ�&"b���H|n�D,�����$$���Ftfj�QW�����Pm��c��#[��?��>��mn���A���*\�M&��U������}�[���RH-�(�4YE+�p�!�C��u��u��;�fD+{����s�9�F{ K�^��\�l��3�S\%'ի6���i���P�I���A1�؃9�ЭE�
�#�j�UQ��$�ª����o���¼ �s���+�j�7&TBQ���L�K@C	�	�!{d½i���q�3]�5�a���#8N#�<�Ml�����,!%�����Lp��)p@۪䪂u�pP��R�v�� ���W7�@�wi�ͮ��3���Ǉ�j�3�nK������î��sǨ<i]gޑU��ڊ�>�a�a�lM��B�؏��N���TMa'7"��~�V���ֆ$Y`n����#LB�\���-z�qc��/_K�8M�0m�׊8�@k@J�\���
[ʘU��O�"���x�!I��[qG�r�K�fp�H�4�^Ѧ2F���#��.�����)�Y
5*[��YGV"Y�*�%��+=U�v�|6�&*�;�l�wx�,_�_#�H����@I�ru�I�)'�%��:}G:/:��v�B~��:f%c��h�c��*g����J�O9�g�lڪh��P0;�}K�s�B����Y�G�k2�_��(5�O
�lV����HpjE��+(��: 0q�Er�7�5��+�9�(�l���(M���:*o�#�-d��4�(h}�J����B��=��y��P�@���R�2���ʩ34�i�׽�Rޜ�9�c'��X���US*�Q)䅞�U��9��i�A�7��'l;Q�߁�S}�����.H��mL��>���_�B �|gV]HѼ��L|�S�ׅ��J�K�U�b� �Sx�-�b�C�y�U��<|��*�A��pvbj�����|ПvN+;â�n%G��X�O�RmXE��r!Q�����`p�6���Ły=�ޘ{͓�mB�P/����oZ�+�G��I{P��5W#J*�ݓ,`����+6\�[OMGo�&;8)�-e�����d��Q|�����4e刻��h�>_�?�1�i��p���/�Z�OĚ���|�u��+i��3�,֤܅H	7ޒ�A� ��^���zM��׾
�R�M_�FkN=� @���l����A ~�0��h:��~�������tv���r#��_�,Ҿ��*R��:W��uMK
���%��x�G>ɤS����8)��=��ɫ9��j$�Fn�M o�Ci�a�)��j	�HU֑�ν0;�v9T�s6Vޢ�Ȇx ˾���viH
l��UP9��R�܊�RR`��EX˙�_VY��)�$�M	�5OA�]"k����q-�Ⱦ� nE*k��J�i�l��C�	�8�sPm�Ω:;~2nY�+¡���h�f�M���n�g㹭����-���|����\_+7�h��yk�U��S��,�`�����~m�j�ץ5�2�'����2��^)�l�RZO3z6@oIC=��{�jhW�'��y�M(���x���z��|"��a�ܔ��#~��4쁪2��L���-��"@l �/&���6pe�'�!K�ǻ.�A5B;:�J4�x��|l���
m�E��j��E�߷������vqNgU�X�zOL�-�=G�u�I}��&����k�z(z���b'XsY�~|X'j�_�Ug�R>��-��ȭu�R�r!�-+��G�g?���9Ҷ���k\��v�~51�3w�Dq˦�
�4&M��ʏ�ǁX/�y8o�KR7n��{n�?���BX�t��y�0�[&��q'_諆Q���IO7�H�Z�F�*֝jU��~��gĈ�PϷk� _�4I��7��:`J�Z� ��Y A�vs�.�q�X�4�{�c�%�3���C���1MI?8���a0����!�]4�]�Fe#��n�%}��7��e{7�����^JOƮK���$Kt����L��S��tDa�$n�F�_���ql��d�<����.=�2� 7ͻ�ߤ@͗' �)1)ͼ`�����sC�d�Ӡ�dyJ(���B/N%�(�8�Ƥ���?td�y�V�q��W�:��g�g���_p$�vꈤ3U��ap�U�f���k�p.�����p"�zŢ6lt|��0b�i����WMߦR������d=��F�)�P�m~b�Rw�-��?�}�u�����5`ms�+>�qRi'�<��8�dBU�/���&�/�E���~����<d�Gk�J�#k��d�;�h�׍�{\��[�v�q��7(.;y�Û�������7���ə� �ðo���^qY�Ϩ+�H�o��Q� �v�m����8��z�7����p?�T����x{�ݏ8v˫t0�W*���CD�k���铟�Ӈ�9L���(fݓ�X�n^y�m�%�@B���>���''A�<G5���Y� �N+��½�i��;�x@�d�p�2�v�ኾZ�ۈ�~(��o_B�������k��6�wޥ�1<^pp�h{B��r�*���W��zV ��wNiP��E�� Fpg[89�Y�����������V�ǷKv���ma�+Ri���y��a^Jy��[l���Թ��α�<�,ۉ*��M~�l0�����"ÝUQ�eB��r�s���"��eUDSu�M#+�ƿ�礶v�c��)��ZY)e�T0�9��������3�gtqt
�¦���cm@֓�)gl����/�V�eIh�N=�M��u� `(�>��Mi�h�DQ�6Z;3��w5u�#eJc2�2����@�� yNuX�?ss�E����vq���q��cdq�}��h̅����C��N�`�v��6EA�=��+���;
,ߩ�E��>�5P�
0=��~#���);Z�y%͗	 �U�o����s�N��B��9d��JW{7\�fT;�^3ظ����H�G3��V�n���8t����ؔd\�g�R��Ǟ!{�P2}GG��3��g!,5�8J�
�.�YϊsHL~&��)���XH6lQ�4�K�������u�`�#R�~�y��\�3��x�M����Hр1P��zorws�v�-㧽U12<ޙϙNr�����N�w�&X|���y�^م0��ݩf��4��1W[�(�pIt�K4P������|���ft,�M�f�+�\�d.�9���nH�I�7`,��,�r��1��={��V f� X��W���g���u������(��U���2�P����p�,��V�,�珜�>��XT�Sb6��}I�Y~{�t��u�i��9|53�o�DY>�hh�Xԏβ.���j�����:^��=x�Cmu,gz�}H.i�*0WK�'Λ/�Q BP��u�ԍ����c���0���W�Z^)>_�,[�h�#Lg�Vt?�����!1�%���d�G��`Ԫ�J䯗<��F����!]�Q�r4�6/�s���eUq�.�K�Qd)G�/�=y���	�#g��:���k'"i<�@u�h8!+06������=�6�3����q�L���t�u����l=����}�>[��{:�K�^�+�d_v��8p#�	d/�� n@Ѥ������{(�_O<C\x�Θ�3��}f)�S.^�3>�i�d���� F���)i�P�C�#����H:
����M���}୅�a1�&���X�ŭ��[��̡4V
J�{̛�*�T�	\aU�G�i�� ��˛��.x����^c W��K�]t��p���./I��7��B��=mUb@��7l�x�]����B�u\i<�ACO4�Y���L�����~�Ŝ�*ّf'Ⱦ ��?+��s4nj�ςY3}���AZv����J�1�x��/�g4H4�%��lx���w�j �,}Y�Z�j0+?ނ���ȝ���N�$$Q����y4�îx�}����Ը�L�����w���u���O�h9�R.�����k�T��_�s� Г�ǟ���&�~U�n�OTe�]�d��ZEG�'���� Ң^;p5��w�\o���m;l\?lL轛�.E�f���!�+*���,�;(.��~�	F��U�R4vgaBC���a*�"�f�2t�>o[�H�=s��"~b\	W��9���y��'�u2醚K�����[�"OQM��	;��w_�ݤ�P��i����Q�5z�.�EUJ=����L�;�\ :��5��G��c4�P/�z�\"j��]���W��B�Ϗ}e*Kp���
�첆��2C�l�Iu������QaH�<�f䵜P��s0�DEYzT��HLI(��J�o�5?H��'[�����[e�"�ؔiw]VNW�[�Ƨ�tL/��n�'x���v}J��(�17g�:OK��ڭ�PPR����>�w��Kmj2���fǯ��"����IH7wz�n����>z�Sg�a��J����.GK%x����Ԩk�'��=�[tEH0�K��J��(F���Mq~��Nz;խ
��c!�lfu����rCl��F�'3�jDt@lL;�,1��6�[QЎ�tk)�iS������p�.yq�8hr��bGcڙ>"$�!Q�R��"z����׏���
�Fͨ׉Ў� M��}�-�Z.'{�-�qm^{`�汸Z&����<�p��||�L�����2�h���|+�[9�+�9:������'Cxq`��1��5~���ꯣ{l?0����V��G5w
�4�6�/!^����E�٫#H��c�V���[�㞡�b|*�_a��֌�TCg�L˺���!�W�Ю��Ƅ4�h�\����@�h�	��??��*^��o��͡�����K��Η���C��5��V�8@��� ��)�]Cm���^�$�F�6	X�~~!{��[	D�&�#��P�m�� �q��=�`Q��w������3��&(%�vh��۳7���,qR�E����?0�۲_KR]�� ��,"�6s��
����0�s�Չ��6J��|ɾ�	����>I#�*^��Ij#��0l��:ח��,8��/����=a�n~q�οo�=� l�#ǁ��T�����2�pl2��%0c����s�0zF�f�
��|\*�@���sUF����#��p c0�M(�5�H�S���<@�?�S,���+Y�B.8o�M��YǞ*���V1x�W����~��p�@�{m�ƽ����HN���+�΅	=d�ɺ
x���N��0�a���2	`�faq�����U���Xg)Dt0J�px�9��z��8�ekӥ)���`d�;���r�ݪ8Rw����m�i����;15@��I\��hݭ`��D���J~���U}A���&��/:ɒ���خ���A�eF�-'ϓ���"P�a��8��
������{���!h����?~����_��t\�q���T��G*������ҩq4�I�!bJ�{锷�C�j&~Q�4t���G�kBz	��m]_�')k��)6g�w:X�l3P��n��yJ�!)�@Es^#���8���CP�L��pH�S�\���R��}����;g�h+2WB�Xi%��/���P��1��S���j��U'���b�pj��A1��}ll�O�vV�S4kw�w
��ذ|����V(�@)�������Β�csB`Q��dc��87���KB�S%�3�6���7p��5��D�ыI3�Wb�2ܗ�*v�:$�lJk�Ua>�t�3F7LL���`wd�ִ����e�=_�5��m���K��6O^0I��dd�=P�7�zx�#����z�L����QQ���d�����"-������tp��L��f�3+�fn�����b��3�q��'g�'�]w�w�,:>&̀gd\2K{;�k|���CD�ذ�jꐝ{�b��lb�b��s���*P	�,����PۻJ���)2��;sc��)q�geZ0�`p�oԽ�G�w(_�&�孥�{�X^n�f��K-�1G��ZfR�l�eT�X�hP7�[�/ ����iE�b���{���Ж�;)�Y�m<���;�RG�������w�QH���J���UD�J�a$�Ζ��o�
B(��[�b]��X��2�9�;IXi�ERD�@4=�*N:^���� �����FoMk���3Q�K�4&ӊN�L��:e2Yz,[�g��t�l5nͰҥgr
9��Q�K7��,F� 4�W����>U@��[v�~�=ߨ$i2`둼�wPK�%����u���HV��kG餼���B�6�9M�$�G�oD(ھ{��"�H�S�7���Z��Q�ӂ�d�U�K��%�����?��2����hv?�۔�X{kg��7Ո�R�� h���k@%�VcL�M�K�(�I�_�b/<���D% i���"%TbAu�,�G��l�?'3�u��g���8XJ=eɷuZ�A����)]�d���X���+u��W<w�(���6H�����}���gH�G���r `Od�HR9Gn�/x��
�5�WU��`HÍ�m��ub��q/����dB��v��폕�e|��4]���Ϭ�2
$
�X����� j��0;��aWf,1s�-��Ԯ9�'�QQ/9�u[Q�rB"ٟ
�z��� �$O��p_%[prMRٕ �
�,ϝ�|�s�Y�^�~
���)�k���u�Lɝ z����} �OE<�C�|I��d6�F>�蠓i�|���K���6e������*�o�A�#_��	>2����)���4�N6E�g����9~	c�����c��w����`��u��2od����� =c�\���팡jI��Bb�$F��eq��M��u�.����ڳ�f�*^��|�-`����h0?��v�\5�����B�]�e���.�^�g �S�<�?w�w��%½`��xJ�OFI����r��5R.�c���'�N��o���Z�k�����!=����̀kX�4��ٺ�Ue�	znµ_�7�:�3dyD���!s� d��`V��^���!����j��ꢷKqx�!�=s�`��+����tp�D�}�x]�J(���E��]��Fฮ�񹟦�s��޹����V�d�bKUw�B�}���U)� �j�?��Źh��6:|6�1�����\���t��DB��!���?[Q�V]��HE6�8Wr��n�Ġ���#�`a�_E-A�"�����X��>(�Q�@�],p���47��C�z���`�_|�o{ڪ�Pñ�e�o� ����)W����=>W�V]�y���lA�ơ�Qo�r�DzV�<Q��4�ɼ7�u�`�]�k�_/�"��3~t����թ��2m�tb+Wp���$��k��94�N��]>��.8mJ���P����4]a��w�R�
�_��`]\�4R�F�~T�СSV}۟��cz�K�2D������Ө�*UP�e�>E+<gp,��L���y�BC��N@\�h�5�Ϳ��1��h�C�����	���=dI����(�
m#��6�Β��D-�1�+�"m?�aLQz%7���9"��?ҵg�|��[�w���2Hj���T�Q�ѹ�,��G'���Q��-����~���J�{��lBr� ��}{�杹~���Ǿ��[A��Q�<���NQ�X�.���R_zyu����P��b�����V�װ�8kz f�C]h>��]J���j���QZ��������N���6��y�ӫ4*W!4[E���^����&��o]֖�?wk��Ѷ�W'������|�U���g��Y�9�n��G��S$*S�k���Ap��Cx��tS���ޑ��S`=��!J�0�=)���:Ki����l�����_��W<��pd@6�KT�O�:�Z+�x��	Q�_���"��jf������XA\.����~�s����2����6�]���n���;�G��0��?h�T>�8l� �M�4��v����������@z�*\��492䬄nj'�R�������`�³xl�M�3�˵�>pa�Re*��I��3�������"n��q/��u�nJ`s�{*G�0�.oӢ/�_*�'"eN�.u�îu�oZ�Z�(D*��q��ʚ��i[����Z�t�^e��@�%~ �hS��a�����8�qo֫6_B�P�W㽖�`Ibw����K�H��s��Z����;ft��/�v}�z_~�+�G��=��&}��Ė�rx��
i�>OH+�>��kNw=S����	?��f�j��]ޙ�t�, �B�.qz������o�ig��K�ք>�ru��M�S�"v�7��:B��An+[.ǋ;��s��)�D{@ז��W��1���O0��^�%�Mm5�^���P]����ʲ��uĝ
�|0����K�o]a�c�/ǆ<w"�B�%��Î�Wꉷ�]Z�w�*/���ǡ�����1���	�T+8�#�P.�\�� ��k��s�x�v��P#D�'�	�,�i�]7Q{���ϓ\%��v=9�|�;2��f�
{]I7̲��զ �ô�!n��5Y}ΖN��>(6,�4��g���wɢ�Q�.��x̃􌶐�����kG����4���d�U4����S=���
uz꽼�Ur���W؜��A�H7�: T������PC<匧�e�'�2(4#_}���2	K�W�-�҅��A���N��@��nā����\����)̓;��r,i|��G�7���!9?F�x����z�/�w��o�BV�x�lz�g� %�A��aNs�y]>tF��M	,����Y�j����!���L��6��U�{�tiC�M����,q�8���c�2yLI0���N��7��M<����zT����/��a}�>�����d�u��a3��L|x=UD	�P�ҧI�w���%x��X���ǯ�?��~����@3���*)R(�Q,t�W����ΥQ����"��4�pa7�p��/�H}
�+]E���=֢�2�Fc/k�.pʒ�S�Ӣ���Z�nj����,
�b꺞�Z����cј�3&��T����>��R��Er��b�B@��5\.c��n�/އI�/)Of�WV�tk[���Ǡ��α%$~$�k@)͖X3k-�1�#
�"[�o�jP�=�9�;�x�󽹺��B�{�IG�}%Q�;V�r��%�yG�gD��l��̕y*�	�t�6һȡ
+�h�T�u�	a��+���D���Ta�3@��6�=e����>�>K�L"[�u}!��לNI$��N0�h��^3�R����O�b�&�a�-I�WC�_?�Z�}�	����B� )E��8����4���'��Ъ,���|��zVTЯ_�r�U B�S�E('�W�d��� @D
�8����A��i����.�d)��]�㠮8�Tceq5<��J���TL*��F.�a�x����ۑ�Np�����s8n��9n�M}k���"�;S0���A�q!x�;w��:�R7
�p�����ؓ�8�k�{��qny�[�j���6g��_p��
$�$�۴��bf����(0!î�2j�8J���^��;�j�E���j;��?��{��,��id`Q �Q��x�N����n�~������B��am��]SU�ĩP��d��R�ȥ����9*�hc@�Wc�x�h���$[�w'��t�ȨP���Oo�;�4Us	�>�3 V�,���_N�v��׫����vs����)�YP�Q�0���G�D�/A��LJ@m� �V��D��$2�Ý|��(y�-�Dzh�����x(6�ޗ���兴8��o��x��Sz^��HFr����Z����-^,Vu���C��w�0�}��?����H��j���`�����M�I^�n.33+T-S2��_�~׵�>�3������a�e�p�!�%���!��=�IR�C�l���2 ��y`��ޝn�l����t�Hw���˓j�z�8;�t�d�l6�	5���@t�0��i�\'��������� ��Nd5�c�%
� ��@iDԊ��m6�uĹ����Z#�S�R��C��|��^��=�6�H<����<�L����A�63�f��Z��3r���y����1�RF�����?�H�6��+<��`�͵�C��o�:���wUHj�O�*���B
H�1���c9i�v�vN�w�(�����&PS:T�����u����o��&�i4XT	��<Z6F�DM�^��1�o^'#D��<H6��H<SՌ���d�]?�5i��T�
� +�O�B��<�$�2l �C%9�:�c�.�X-Y��2|]���JҘ}�Xh$(�C�n4 ���ݞ6y�i����*��Gq�jwt�ZU������w�T}0N�%�'�V>�
��@�B��>J�K��xÇ�^,�$�`���5�C�c�s+4]6V9�J�h��aڐ�X���ؐZ�'�`�9��k�{��]�����m�k#��p	��GNڑ�5�>���@ф��`S�k��<��y�w��x��K����ށ��5b��z��(�4 ���K4혥����Ԫ�V6��@���`5��
C���uq�r%2�Q��1vfH
�W�Pz�^rELp�hF� 2
�JEaQp�bd�66�ĥó�X~A�O����[X
��KsHnqA��+L`4�C��x`X�������6�� �~+d^�5�m��v��iauj��LN&!�ɉ�*W���ه����ԡ��݌���:����:pGW�Z�[-�Բ����g��]o +2�a��9�&[m�0_^<��p�o��$2��۬�9�6jw���l�H���ol<�LCzr2�@����K/��f_���'�罓�pQ7�T1���x���������>[Q˹''g�]g��|����{!3��[% �Ț&
;�HdQ�/�o|��a�L��1�]ɗ�W{�V�I��B��lS��<���a�(�%? $.���m&�e�-嘥��U Ğ�_/xd�ϗ+��^��l~�w��
���k��Ӏ>�5����J~���Y��+�jQ�}�ō�oI�FSD���q�|{ހ$1��� ��*\�wY9U��J#�v�tv:�m��J:��W#��Ў�����ԕt�/F�
�y�J��Z=��䵅�蜿�1|`��u��'!�.�xv������B6����j�e���i���("���K�,Ԫ+-A~e�ڳ����0�� Y�mV�<w
6���1��\c�( ,nwؠ�=vm�PԿ�Z�0�<��8�n]���K��Os�	�Km�'�Ŀ��/�u]�����}��?�$��<�~XsIO�n^�����(k�M��r�l����=�cK�K�yik�ú志������!o�g�2t�z��/�u(�tw��
6Z��"�Q�:u����
=}Y��gI�}
��.8���(�E�lj^�h�u���X�H��G�я�ŋ��o����V�EG��#�!x�6 ������ <���m�2����p �U��@�ޫIK4��(�ؠl�Z�S'%]�F;��/��Q�K=�]h��9���m�m���C�z	�����7y� �5H�Ĥ˿~��{�xC��9���� )� ��N.C�ʯ>��Jm����~x;��&T*��;�U��6��F}�Id��F�N�շS�p*L6�l������Z��'��rhmaF�5)x�����S�=���̳�*�t��O��+�%bZ�x���R/�	wMRV�E��O���qF��T���F��K_ł��44گ����3r�k��ߣE�"5I-��An��D��?�����V�B��qPs�����m�T��#P��Ck0Ho�p,S�m���4�Z�aW�,����(��7I��_w��P�!k&�C��Q�d0w�u_Ш���;Fܳ���0��μۇ����"s����A�ai^�Z��4\���}v�19��g��1��B5�o�{�W��&w9�֛^�f�Ů�P��N�*�9�E���]�s���y�65�I�a�|�����$��*����v�D�^[�-�}�[�t�e�ı�~!�}g�,5����eM��?E���r�1"ƹ��k�a�\p�y%M�(�N�]I�^<�5��tW��7��c��]癔�]Z��T6��T?�_d
7�#�v��/	G��d�
��2����	P$|{G`��Ab�d�����;翌��0�X��pZ��%�-�o�#oϱ�\uJ����7YUƤ���Y��sc_FS���9Km'1�g�3��hk����G8�1�\����~m�b�&>p0˟p��5Io���aQO��R�<��̖끐�Gũ�u��WyZq�^%2u��|w" �ӌ�g��������R=���d��&��+L�=dn��F��GV��q��yK߭�"Ӵ&�:���L��O�P�#��z��`= [3��筘A~�������8�j���V0	�	;/R7谵���|D����aVFa�id���~�q����\K�C���_%���Ҕغ��i���k�z�`!A/z�xbE�p���cϩ�C(g�-� Gw+^"x�󑞌�Z�"꿝d�d���Q�Pp����h#3���E�ߑ��N�=�f����,6=�$�D��3i(~E^��"b�I����p�_��H7:�2.��,UTY�a��'�.N��A�޳V��eI���Tذ��=9�c�f�|%i���6Ͷ{�ЧF�VW����~_��P��~�]OL�I�L��`���������,����3���g�c ���<9f����O�P��y%Nix�G-9�Ҵ�i���XFG�n�F�`��w��pS8�>���k%�զ��[�B!­-�3H��k%�/q�5��@EM��w�s[�yK�aEzEQR�u�}�Z���{�zd�Ѯ0QX��Ld�t���~�=s�i�dd�jc'7YK)\�fI��љ�2[�{��ʲTdz�x���H���m���MahJ�_���2�қb�:K��Tclʼ��	�gZU{l���ޚ�ek���w�y��33k3�<?T.�w{�c��)AQ7�`<�uC��E�TG^)O��P���p�w&� ��I�4��#J-����܈3����Y�A`y����/ؗA��8c���\��qR�S��; ~s^X����Uə��N�E�I:�;+ Q�܊�������҅��3��;��a2�����G6�tf��dnC��)�؄��a|��W0�m��%w�s���eH0�E8*:"����b�zr�9�f�M�{ Y��!�;[��5*�f΂�j�Ͻ�;j~��"���vY_紝�>!���?9��M������"�`g��Ց�^}�H���'��F3�A����0��!�ɹ�P*BV�SA[<�$���kY�O�4�]����~}�<'������ƣ34W��̅�ef>�}V&�? ����\Mb����[�< �ƀ�☵	�4n���sq�Μ��+�X^^�i&*j�'��F�B�b�FP
���?���y��t��%�i?%���r�I�C1P���M�B>��ᖇ@l�p��ѓ��%�5�+�?�<z[���M�����*��j���ۀ#SSU+:��%DUBN�� �|�S���R;��C����R�b�'/E�}���䄄"k�h�m4��C�|��~;O��hl��u�C��I�����0x���H�O�g����T	b0��:-#G�5�:�|+8��(IRo���Dz^^ـ�$�%GK�&~l���q3a2E��6c`<{�Z(��%�hM;�+�9
��Rʴ���F.���hd���O�i�ф�͒����L�h�� F�9����00>���~3�>,AlT���S-�h,�4�k���v��?%1�ė�3��Ni���z�W��D���d�<�������q���'�Jw�k$3������Ńԅ�V]�yRpF�?�� �z� ڬۡ9/��sAEN�Κ�de�'���)0��I0csZ.a��s4�Dw��XlyAW*��kb\F�t0�D��ZjZ7 Pi]|u��)��GvIn4jK���j���YΡ.Ɨ��O�#u[)*)�=��v�"��@�P�Ԙ���F��V��)q��b�rخ+e��_`�9\��=�8N��9�h��q�tq�v��b�kC���Z@����v�K�??�c���wK�s��:G$ڵ�(�Q3h�s��2�l��-��������0�[��l��q�}'�C���_�+���޲;ؙ�;�;ש��!Q��=Afu�l�pK���9�zT"���	dw�g'�[X�c]+@�����#�� tˆ��=ҁ���j�w�W���/.0]X�k8>d"`8}a��l!�
�����DBљ�#���p�\��I$2:W���q@Ҿ��ͼ#���	��db|V�bBD� �� ��K������,�7�{�Wj
N��]���1�D��CS������G�{4p����vͨu"q>V��������V��'�Q�O���[���@���]8���Ǟ4�K�"{U����"1���v�pX��	�'�?�ϊ��XI��o�bwO�Y��O�/(��������7���NtZn��H_h�w�(°��nQ��f�{��Ҥs�t���>��k��9 ^���/p�9�8c:g�gwtr�_W��-�qWڨ��_n�Xu���e�X6`��f���ޠ/��Ex��B�6���y$��߃�fJ���FRw���eM�_��V*Q���}�M#g����{=MQ�T�&��� ������0�������db��t�0i�
3�šo�?�������Lm#;���i�.t�Sb#��)��uV���B���M�C�5,���_���z�5�2q�z�L�����wK�~\��G�⠣�x`����@��h����s����"�Y���)������+v:������{����l��i�݆�54Y�gx�
[��I(�TJ��?�z���o��׻W�у��0\]��t?ti�`���e���^\"f6C����A/v�����������x�s-ɛT迈,v	mF88�A����(�)�[�Lw�nf����8f?ܷ<���'���0��͓���LI����k��r�E"����L|��Ȼ8��&T<�l��,���`$^o�ǺDMI��{�u.�����6�
&���s<�%i!��Ư���*w)�?�!�ǃ��'��+��e�W�!T0z�gɩm ��H�vP6=�4��uE�Y�i@e��$�*=-Ai.�i6������B��U��W��{��ߡ���w/8���i��_F��<�oM-_~؁%�]6?����W=o�f�{d�l���eܽ��yyN�$c��]���(���~�#*I�Ko�5ND��2��w�IWc�|�����0�q)���H��
n����GlڥӰ�yq^�V�m!���$7�1��J���|���ķ���:%<�k*u��i}b6�1D�����Eɭ0_T�d���?Mlr���gB�ˏϺ_�
������KLBB{��eH���x����"�TeS��HȀn)?N�,�~��Z}��b���r��#�����~�jI�3�=����N�T�H�AҚ��0��ҙ����W�OhֹY��N�}�4 O�wзQ�]����_�$K��VpW���!P���S9�����M�꙼��P�@��� ����28� E�U޻Y�-Dd�ې�8��c�1�M�QN��0�p7��E	��j���x�1���h2�⽒�!v���1/��ұE��K�g�{���ddV<+����6���{�S"p,�zDo�9�*�TF�pf���)M"�(�����D��s|���@�;�0pL̺��Os�˯h�䄚�&��yO��[3V�����*vش�����`|���`m���@��4�1�`���1U��x�+j����UR;�55����܉�5I�%��\�$�<���_~��1��K��k$�0�Z�;�ؽu^d��j�\{A٠���j��B6��%b}���?����ܖ}=>�M<��kBwKy��cJlrUً~Î�w���?�]�W�j0����k��`K��ԩ�_��
!���_��q��hh\)�R�x�C��d*0�#c�O6��1�7�:5��վ���B����<.�b���y��MA��c����D��X=}k�)Zg�� ���x�aM�v�	�'��Y>�ߐx��I򙲃
��dfM�!��s�"wt�����,�Eb�t�,Q�uU�I	o۸9*�]������@�{"��F�-l�_gs�Aᅛp_�|�z��(�,Fщɾ2�� H�k�?���.Ϛ�Ȭ�\�M�oV=���4=��b��9�c���w���/(E�����7�O,t�6m�!�F��`ۤ4	�m2�n�T��b���Lw��u@SL�{�d٣��ݹI��>�;!�YD������p�ߓy���dT���2z�]�p�?j�`Ή(�"�B�:4�֤W,�Ol�n��Y�S�5����KՄ��h��������K�#�xDj�����C9Ԥ�o7��Tj��-e��ީU
��Y��3��R6_�?�(��m�� �g�c}vx:|�M��7��F�*'O/e`�j�
��8(����
weŉ	=B�`���!�]����cY��P�|���孱�ӝ`v}��pj(W.q�67B{W�
�*Xr"O�Q�W�jD�o>ۛx�&+�'e\�	� q�Q�f>`��8{D,�2�<l���O���b)h��_��_�����rz�^[$D�-J���Iv ��!_}��NO H����X�ѐ����Wl�n��V��q�m-@�Y}~��Ԩ���rZ�����^�:qK�}+G7��(1���g��ΐ���dD���-���"F�+X�]}ѱ^�S=v�&`dsԓ���'�^��A�o��|lg]���C.��jpZ�߲GgT��߷M�I�mJ#�򵕃#*R�V�'"D6�� �T�J55�>#�49{] �*h�z���/�^�k����x�����T����ϦƏ}���4��2���]���&��.q��t8Ώ%�������T�Y%���"��u��${HR�g;	��W�H^��8�V��֩%��,Q�vx0���g(߼�	mj HO�R����K��t$���=�8��cL�n��(��<�~d��~}�8ŁӘ��}��ś'lS_q������7�S�b�oxd��&(���j|�\�޻q���܍8�{�%}�/�2e"��\j�Ol��S �_��?�D�1�rD�5�O����匯̗o���,Ƣ�(����Z"�.b����OS\r�A��sАl \4�0�� ����r@����d�_�m��S:%Y�ٸ���%���H���#e�b a�b��=�p����嗵�|��p�%�mT�Ѣ^� �%$búV �n��C3��q��F���nm�NτZ(�R+zn����)W�������2��)���t�h{@���.U�ݣ�=�[
�}�hL�e�Ϟ�)%�Q�%�8�Zj����!�ۣg��˰����	��"����r У��(��[:G��<�i%�/��*��Ԓq����4C���A�]����q��'Z��A���d;9�ʑ�Á�|�`L��P̻F�찝��p
x��W=Dw�����Z�it%[��ؘz&��0}DW���8�ޥ��,JK6��q�ra�k���(;{)@г=��?=�K�C���g��{���b��Y���A�'�Us�O��ꇨ�Dy�q� =mo�r�����/������|��/n���_�$�*L��AlHw�d�|����8��ݮ-Zm7�/���Ĳ�	Ld�T��ᬗ0��#�Ѫ�-7v+a~�F��'�.d�X[�I���5渝��$>��3�v��%�����0�?淉3 �v됆4'r*���7��kn@2��t���&[��F�nm7�-��q���!zw�Ul�>��) �fs8�T��*:s8��������{X�Xؖ��8��L�f�G��C=/=#���<��q�_����Cj�=��
��m+�1�X�e�O�� \1�b��[��V�����Ӎ�xp��@�eͨ?f�q�I�{��zP|���� v��L�������dۼ��a�L\g��֍��^gyR\�p[![ʄl� ���T�U�c�aJ^���þ�kD�,_��$�l�d�<NYTv<�7���.�&�pa]���1�ӊ�1ҩj&+����؅S���>���ք��Tz����Ǟ�8���B��0��pcA����LXi���ރs]�L�&3E���N.���4R���S�ad�홚(־|���`X?h<��1$���j�����W^�7ڥ� �y~�0���a�C,怷����AO��1J$*k��akDR9�r����|�������Ki]��6��<�"gQk���uH�/��1jT�����3'�`�/�3��[z]3��5�e�r#��)e(!'��v�'4���,Y5�Ȋ�E�8����%dG��n���>|JQ 7	���hswT ޅĆ�+�nK�Z5�$B���u��u���3z&�V�r&���GH#)+.="�3�D����'�	B�E����&���C���ǾY���� ��>��ng�Lp�_��E�����L�?�&�_��o�c$�0x�g���A¤�}�r��������S�B�ɗ	����S#~�O��=�Hk=�_ �`�"꧚e���~�2��t|��_g,�g�����?^מ�/� �!�#�S,g�3���@G{��-ރO�w,iwhc\״���^
����"�R��"�>ƾ���w�xqsB�J����tY2�qB�4@���IB'�i��H<�db�b�a �מ6�1<���s�[��XN�@ZDUy��d`θ�1C�� ��RB} �(�|���~Dݼ����#�~���&������,���N�f\����wz�9.Doh��d-�r�a('6"'v�w^�����Uz��r�5E)�������������lFr�}�@�',O���K�G�������~�����{�͹Y��ѫ���A/*��w�ꁛ^�[g�m5�N^�GܖϮZ����(�诡���ozqʿv�ݻp�����8U��i�)Fo*H��b�S��/���:��q�K�p�b)�q�+OL%�'�FIZ���߼y+j�T_�M!�@u������g��ߓD|��<ӹL�a6�~�(�S���ZIr�_?YN��' ��+��,Z!���ՙ	�0����*їwP�����5T�%L��ɮtI���㬾"?Fsu���"ETR#<,��.J.���,�m�!�m��P�4��G
�k.+,F�p��`j���-4��"�q���`��r++\��G�h�UW^r"�$���N�[��/@�:�g���eԀS7s����k��!���|<n}��d�� ����s*��~k���Yъ�O	��
<�x!�F�	������&��1�TQH���˪�L�r�x�>�/���}v��4�Q�Q���#1D��ź���?9�_�H2�^�IL �n��|�BP0�7��O8�%L�'��DRH��>3juB��j;d�P�����PG;�Հ�S�چp�|o�
wV��H�8��31���+���:�Ͻ}(�kHN�13az�hF��{�%�F�0�v\�$nB<����3�����0��9��G�'��������{}�9붶��L������:s[BbV)��
i�Y�,N�D�-�� �Au +9�Zr+vf9{?�g2^�z�_&��!��lL��ꝩ�>+Gط��kOh}��d�Ӏ/�c.:k�qf��Z�L��oth������ �g�GB*��r�)H�Nsnz��!Ns�?��K��k�`��}�
!�}F���㚜�`�S���E�[���|��?}��;,��u^�P�ז!3b���g�2��e%�P߿ǧ�x�5pq����<�M��Vt�p��<睮r�
��\������cV��a�h*e�8����BA���������0ԅ���^EJ��^�Q�ƞh��$-E�)w����/�&r�k��Uf_�x3˶#��; �p �-�HX2�ȠW�qK�O�+��o����d9�@�$�p-g$� m�p�B[C�~�?�]��"��-u��B�p�Q�������Ω6R�y���t̬>9��Z��dKY���?��t���3 �)5�����[Iw��T�	�i�04�J��SC���$�U��{s&8�	9Vb�N��?
`�N�z�?�n�t;��
X:�:����S��z��])a���wu���
%�>�$�b[�1ш�I�]�#�D��sy|�g��j������nޜ���g�U즕��5��o���C��j_PI�T���IqJ4�Nŵ�k(
���0�k9�$$6��[-� ��g���C��SB�/A�����ϳ�9�/_[rg�'��<�07.�o�������d��ĥ�!V�{E�B���v��AKIkR����v1�~�vvt�w������Bt��q����7F��
k��ُk����EF�̽�� *#jN��7�ǰ�}8<�d~��[���s=���H)���]��g�S��-j4O���
>鮷j国����z��x4ZL���|A��0Ϊk�y�
���ױ����\,��1@�||J�����ti�n�#��^�T�XS�Ֆ���43'����XZ���[��6N��q�nc�}쥎�V��"$%�q�V��G���E����u����y���l`�|>���6�X�#F�h���6z�\Ly~�f���t��[���5�«���\ߎ��L��=#�U-m�8��t�<"��&�`�~O�4F4����#Ø�������Ԩ9����~��%z��+@=��ԗ!k� D$�Tz�W<9l�9^ �����_���<����`��|Jo4u���B�vL����:����?���|�V�`^.I���3��� ���<G[s��`8��/#���WL)�A7Gkz�Lp+ѻ�3V�b�g�7��뷍�� )�����AZn��a@��r��v�*�YHSCKb���R�6g�y��hz	M�ŽXB%�å�B�k�U��M��1�>�a }�ڻ?�2pt�kO05 ^��P7�%S�?(B%_�SU#��	�:`S���R$NE�.�M����%O���[����-E�/�hNn��u �[h3��{|nY��ɫ}����W���.O4��<{���#���Lzis�I?�4H)�.�&�$N*;�?ޘ'cK_r�V�{F�G���� ��a"��KYT3��d�X�Y�Ak�����No�
�`���IC��<��� y,�}!N	d�_!8��Tqx뇹��v.�}P���1'X`��MI��z�F��kO���郛�o����<��_ҁ����jSB�|���Ea����]%����.wR�^�[ �NP�id#�t⒘�{�_>��0�<c��[����{�ʐ�?����:�Y��19�u�l�=�h&���R�t(Cs!(@y]~h�d��!�Eg2+����y~��¸!ԗ�i����Mp�m��ܞ���ՂH�3�����:�hL��'6K���	���`�_|֘�e�������&K�E� 㷓�=�f7P��P�)��"��(m��2��r�Vy�}��/[��zx�@aR�����{}N:q�y�nV���&$B�^ǌ�񕆒2�	|ŀ�n{�}LX�r2�`�|�O4ƥ��G�}��f�{�V\�5�Ic�>&�֑~˯�ԣ�,C$�/��	ɨ *zt0��K��Emڏn��1T.�殻Z�|�_B:�ýIR���s/�ȐU�G( ����2G��G˪k�Řgl��Cgf�޷]�����١�����읶?~t%C���͂?<��� f�}W��8-P��Oa�h��uuk�=�FcC$��Q �6~x7PU���휧o�݀���z_6��*�X�`�;F�1�^�ï�?��z�S�>6����0ѓ����G�ط�j�8u�8;Ca�¾8`՛D*顗�S=X��˒��^��a����o/��Y�+��F�JN�h�[W�S���8X�?!��P�Ni ���#��C��3?8bZ�rp�$�J8��b���A�-�Djӱk0]83\4$�"WvO���[��&�/zKݼ@4�wY����5�V%��=�,���B�}�oj���RE���y��q�6�S5�I�pa[|2<��-3I�L���SL���w0[+Gs�c��3H���܁��g���`*���4�`Xw��8��1��q[#�w,e��<-[\s��ܧ����j��0ur3-L�����-u��wׂ+��=��,t�ƶ����J��N}�y�#wH=��\���'`䅆�F�;��\��ھ���I2`�$�!�d���wM�	&� S��>E+՞�1�±���
�����]��W��!�����@<��$U���0�J���#��{e���a�S��9��(�aaxÐ�k~�z-'�h2����{S���h����ٓ&X��+�� h3LJߠ#�e�����u�tS|u&�_�;b�Ǣ_�,(/���?�������/\�!�)�|�b(߾�s��Z��ņ�*["^(]L�z��#~�adh�vֹ5ڭ4���e�����-@�e�(ٕ�Oq����5P����O�Q�y}���݀A0 $��T�	�s�2���J�cH���vV�Ҁ]9j^�E��d�Fg�U"��=���`�I>,��p����<SK�;v
$ݠp��#F�.*�)>�퇂������*jCR�H2�����=�����@�{���:�n�6}�|�I�D�ݬ��FMz����$�_�Ά�k˲0��c�:Fxs�1���}5��?�֢�S�x4Ѐ�-�&W�R���V���]��y�e^Ek��N�WIٍ	X�|�}����K�`j�Ҹ�b��`�B�� �'�[8s���v.?���5#�Pr�m׌U�'���z�F���֙� �����אN�QߔQy�g���m�9e�#�\�lu��=���l�MX��q��2z�b��3�S�B ���#���lx�(`�3��%l�>�΃�@������!�2��W����e����7��<��,,v��9
(Z� .�`�Yr7�m�a��]]�$�޻���/ҍ����9��H,z���"%�R�a�͒0���_a<�֗{�xʶ�F�b�fsn��/����}Ũ�D�C��q���lKC���ĭ[�?��CJ��N6t�.t+��	/�ct�0���4}��Eso��7�#s��46�b�bE���������k�ƿL��6� ��@.ڨĢ�x��j!\������|&�X�`�tǢ���lܠ6�%�"�Y�C��(:�r�^���,2�׮]�]x�������=fl�O�
�Ci���]��MY��SF�����w̲-�o
5~�WY�Ք��\&�9���Fõh����&��:� �"���
�z������Jv��{G}��9m�%���Hz)L-�{�MZ�y�[��d��X� W���b6��A�ΡS%���t@��Ɏ��鞧8�NE��@�8߲js� #��Zi>�S��nx��� ��a��2I_�y�i�g�W#�x�&&���@�!����w�������%�V-� wT�?~Ҧ����H��^Z��Of����9����i�?�lBјj�l�e�?n����fI��;s}�q-�[ד��3�f��C��^��,U"����FBr�!&���H� �7\tf��SE��F�9�t�~�V��
g�t�cMG����	:R [�����7�;�[�H�|�Z2K�@�[�yLpQ���v{M� �W	�[K��!�V�v	W��y�ס�����D�t��5�,U5� ��Ǯ.��-{�xH�H�[����D���(�>ʡ�O�DP6h$���u�ah����]f;;�7?ӫ����:�}+v�U#,a��mV���3;|��<5�,tNX���(1~�E�G�=��1�i����e���H���y�&3�P���X��v����"4!��N�����DG�1�����SQ&9Y�r����X�TgК�^���U�ڒRN��$��Ϝ!�)=���$8��m��gԜW��Z !���l��c[��0� d���c��1q9��5A����c�6]�6�d8{S�2��)�1�u�!�m]^<7a�x &��0ɥ������dW �k x�k�t	�9����p8N�#/M��Ԩ5a���oZ��q����̎ˤe&(� 6��˫���q�W8�M����s�a�	� ���ތ��?���;��0w���3��**��TD����O�G��2i��=u�),��Fd+
�L�h����&8ڽ����q�n�\Y��R;?����ӽ �`���@��ۿ�[� ���3p�@��ʹ~����K?�	������|��bY����w��Vť�����0����U��U��7N�Ő��jE�`�+Obu0*N2���P=�$Gc �Ѓ�I���~kpBg��P��3;�ٯ��	�'�a[�����ҷ4�������b1�¾��o��+�Bf��$T���v2ZX�S�����sS�u*ެ�k/Uk�*�P�(�ːN`�R��x}��9	T����p�Q�΢�u�B���St�ɃHF�eek{<v�������؞�5�Y�e��؄�W%{�ye��.���h�g�x゚#�����l�H�����=�/#�@|� ���|��mJ����O~�#�D6G�7΄�,�%�D���y����E��� �Jc�	@����m����,������z��>�ȉ�L���b��w���M�lu �$�TM��yT�L$�{<�iwެ�����~��Qz�u�~?����
�[+�=� ��U(/����i�!GTo�+'j�7�ag2r�����a�eF�!i�\�{v�7��F|��u	��^�T�1-gS�i$�j�g�p����i l|�pR
��4��7LR�
��Y4V�Z�I[��'fG�^p��F�r�Z���U�eⲭ\<�	�X��j�����?u;���y
m`��A2��M������,$\Jِ�x�>�է���.�A�bu*����K��b {���b���{�m�JɊ3S�o�m��j��w`Gu)*�$%���ʼ]
�����Y�T���<=5Xwq -���m4����h�˖H�j ����L/�(ӿd��22��0�2�P\}l=l����j�4z�����B�_-��j��y\ �Cz�r�8�\�1���O�_����������6'[�*PZ��<9�����7t���O��9Z}^�q@c��|Գ���|<�mRM��+"ҳE���JN��W��j^����`��%�9����Dq�xl�o	�y�>�o~O�>��UC�]���'e�~�l�"%�'�($�PNް���Q���)�i\����F��m�˘��S}�0ɭ��<��SЇ�}t�
o���7� ��7�%k��g��ȴج��0Z�kZh;�T	�J��y�(�Y/�w����XNrLն��:-�A��1!�n��WH�?��\P̉q���\(��!���m�Go���SM��?c���ϐJwՅX�ˢ7X�`綁��m@Y���y)�wV��&���RZ�5u��hɑ-̷;����S�v���nS��a�(@v��_��a�O;��h�ƶ��َ��̑j�z͌�B�#GA��3�H���ʄt�ܬ�D?�)Q�A�L�HS�/���nLG��S�kV� ��J��f��e��c@{�]�D�e#ɐ�k�RV�*?��q����-�;'�Rϥ�5�瑐�Nk�l ��FW��;�v��8�Տޗ���W�RB�j�*y}r£G!���hݶ
I�6b�IB�(��K�Ǉ�u���f�#��hXk"��`f�n�}>����M�j��ua�T. q�0˧���*r��DND
��(2�>9�t�0w�Q�݅I�}�J�P|�9e��jV�=IP���p��?�������Z�7��j�@5������cc��O���%���Q�Ub�_�Aq����5G�w�dp�&1;��-+x�K����ߢ�����|b�@�|��bk���Ӛ(�	�,���(0�� �Ff45�}�(RFJ7A��e@��1a�c��������Le���y������@H[����:�3an����:@:	=2���4>�ؑ '�WJ~�O��E/~�݆����hiH3�ߪ�t����>�淹8�xK�`����s��reh*����fp��j�J����.1���|6�|֝�0�0�����PҝˇH�{ �$��P���
�8���Z3���LPEQd��R�ʊxԉ�����q�!Պ�"�ֹ��0W���+qQn#���L�H�xכ��1yV�@w2Yzŕȓ���_Fs�4��18���:��4l�+6>e��tHc��&ك�ۯ���+��(A�;[{N�*�ؖ����+�HP������v����~{�e�tEJ4;��s�Ip&N�R��}��Z�5�ov[8����@�'h��s���T�:��u����_D��u��R�װ�lw|7i1�6X��������.��Ԋ{?��hY(�m	�昹�5L��T���;�'�dpȄ�"�n^�Q��z㟙y��x����3����\��Ǎ����${��0@M�dj��f�)x�.n�wK1�n	�E*Q5��j�Àϥ�PS}'���OSjd���ٽ������͝��#��Ռ�O�ƌ0ی[<ȻXd�)���rk6���5��E_�s׉��9�лNm=�~7$�z�թ�����q��jI1��>X�����~��c���.*�:��q�y O�Ě�l=�Y��%�5$�=�̔��I)�JQ��
Iꚪh&�B�ʼ���n�k%��!�7���6[FP�mP�]��AT�����[3H����t�#HcP6�����n�.�>/�	\����u;�LI?]Ă3!Q���`�ὔ86��U ���vdE��n[=�;D�
��w�����N퉺τR�	r�r���|�U��_��ւ&h8=ĥ߯�:ۗ�փ�H�{�F��G�Vf+a������s���؍��s	QI��������Zj������ml�Z
l�b|W1�?i�+x�NH#�]+Ie�!����$n�G7�Z�m_�I���6�qY���K��H!�x"ͨ�y�m%�'p����	p����5���b�W�0�a�Ѧ��@��FWV��K�n	
ۧOF� O�\���6���Y���ihfA�)��(�~M3��zrW!<��*Q�P�A�����V�W?j�`g����D�zʯ}>U��*?�F����A�erFw�@�
�K,�TQ`�P�}����)����A��^};��@��Z�j���=H�����Ql&�0����PA���:K��c_��i'L��ZbV`�u�7B�퇙,l~�k����h���ʹ��xE���>�K��9�'�)���t�kVK(��P�3.���]{eB�4|sg'0 ��CN�@+�������M �����x+&Y#�Ȓ*��?���[�D���K���U���"�*��yᱶ�m�"?�jf��2�v���Q����4�F!Nt�հe�0�k،GX�]���]ŃM���"�p���!�4�� Ih*R	����LD�]�h`쉤&E{�8��-�!�4�꼑��mn�6�J�d���9��L�8�6k�ŭ,����]�8�=#4i0�j�k"�]�P����������l�"�ԛ|�;��%Ǳ��\M`a&����2�0C�z�6����'n"v�:)� tz�	�Lzv�"�ju�&�p!�'o,9�\�;l�8O����. i�ߡsQ�x�ecH��1��?�ڸA7�?E?`S�_�N@��������>1��� a���'�P��L�;�v��ݙ����o�10G�n���%�)pBƔ���xK�DTg���K�'�$�,�m"�Ә�p��[�S��t��H֑[�=rS_��h��8�}|rՈݕv,j��P����MG���� J�L��P��[�
4z��Cұe��3Ĥ�����v޶n^�2p�Ϊ�Aii_f���|/*�z�S~ ��ESۃ�M_�/�Ո�n�w�=qA|(�%�W�=�G\�J����j�>��#ۘF�Je{V�������%-��j��$MO��5(�����^=���!5[�����RF�vjG��?���$jl����q�']�:�vD��x���=_n�[{	:q}��G�Z@����mK�H��A�)*ƆW�@�����V�&�&�����X+KL}�#I��b�����6�Y�m�̓ChԨ@���S���w�/	>����}�=M1*�A���?�`|�����K�NZ4$M�'�� ��m[��B������d�-,��G='Q�,hs��W8�"�����Y:5C�%��=�QK��P҇twD4���E�9��p�/]J���u��i�>D��P(L�A�n
&7�^=���@�Z��790�Z�ن�31qbIβc����\Ng@�������8vD�$�����m���\.���DQ���=�K���ԟ�(G�3�C�.fdǻ���;q���Jg,"�ٓ�Ex� u�`���u��VU��l�o� w�'�v�W���'�%@�H�#�HCHP���5��W���qezq�����M�"'w���A�����	���%���tKV�g�͜���ɧ&��͐Q�=�}<�ɥi�����l�1�D�J�=H�t�6�=%�`�*� ��a�Sc�݋Z�#PgX���6�x-Z�YU�"]����܋J]���X�3a����PGvӌ@�Oq���6��+r�a�yl��ө�2e�L��I���8ږ��Jy�K�����'KK�� bÏ������6ʱ���Z��e���(�w�A�3�9t����9`y�A�y��?�|6�MN�(&@5�Rď��[1q��#r��g+>KTz-��J�?��%�������,W~��w,6�M�M�L-i��݃����5�@��v�´s:~?u�rr"(����~X�U��\�yC%!�kx�l����wT�o��I���E/�~�;R&�y�Jn%�yr2x�)]Uc�lt����@<��j�;D/����IN�h?������1��ge`C���A��uU�%2]�)�����d���2>�
^[7���k.�Wd2+���U�����EQI����Z�󳄧��l�0�C��SaH"Lq�,c������eQ���_�C7t�I��B�鄩(��=�B3�^e�
�G��.����N>����t������}��E��m���=�^�BT������]+�}~l��q�<Z�U����
�;ԯk2Z&b��1.���"��&�Q�w���Q�rԕSo����_�굿�7B��υ��W@y=�j����|�GتA�$�U��q����eyr
��?~H��U� ��Ov�K��/�I��A��æ4��P����V6�'�ݤI0O|�Bx�ɬ����eh��.m�!��-�߅%m֝���O�x���m���*�,~�̕ 8�	5+o���lr����b1�Ap���kt�(9c��$��6X�4b��^�1ޟ�k�D��8�&������g��.ա0�.�)A
��+���M9ZKwJO>gL�����T��ى]��ܷF��<����Ґ�c�}���-1\2�����-�E�\HK��2�f�ٟ��vB�9�
���c�;P���fU?i�>��w���N�7�����.��ך����+7�)[��	�!u�?�ȃ�flt��
~�W��4.�}M��L�dY��䐫��t?�]^�\�]F��~�"���
>���p��_k~%_�r����7�IŁ���м^�8�Ѻ�[e�l����m���|�I��UH��� ߝy4�A4cM���g\fZ���uT����z�m�:����ُ{	;�Ũ�/ ;-|*�qo�9v퀍l�?�kǒ%U���6���x�ۜ�*G��| ���ւ<�:l)�8�j�`����� ;vY?�G~�ޑQ�$���3��^#�1���o�|_��BY��%���1Jޖ��^G��0�Hw�1c�+�@�lk�6�>�&�2�N�!�>�w���K��a����aU��_�*l8�Tϝ���&ʓ�����r�> +��"��{����u���RѤoV�J�����G[�&L�"�mc,e/4��M�A0��4�Q��s���.�v�8��+pmF�GH��TZZ�J��f%���Ԡn`麗�ɟuJ/����o��?�����Ңj���o�T���Z��˶+�Q������<�dnˊ�������B������Rދ!Pj���K1��r
,4M��"���L2��T8"Լ$��&��"�5�R��"s�&ZP�I)ZZqg g#F�����Ң�/bO����5��$z�3��� ~��k5�A������?�"T�+c����y�|/N(Hcl�߉�� x�_ZT�gԌ��=!Z�s���׸��[��+�,���w�y���x5Ȏ�f���V?Z#2�L�s�����C3�g�����[��xt� 9F���'�POL>��_&����Vv#o��g�Х�X -�η�?���߇sA��j�x$.d��u�Lg�κ}�g�����㥍G��n�z �Ü�6`z�m(䫺OCjI�5�S q�Ɛ�Clΐ�	��V|��YI_�гp���(��|����o�g�������������H(��ړ�ʖ���ԓ�K8��+��[,������B�Fㇻs���d�yxd������E!a
�1c�靑�z4�&�����n�^6P�����הH�9����dp�S���o�"E���ě�l��\�cn�Di�u��.��0��0Xz�~�6�2��埯;}���ڵ""S읭<��z�pAO�k	׮9a�K�פl(}��N�}�l�9���>p~o4IP����W�d/.��]���^~>�*�CA_nҰ�mOw(8L]�-�M��Sk�l_�	U����E�8:�'�/�[���/�#@������dI�̖�G1�;�K�D���v��A�Q�b	��<aߩ	�g�����?%ȶ��:`��R�]~W��d��;�{�����.�v�*4���)�A�r�@P���<��f�xgC���~��e�9��׫0��Tp�A�Ȑ_�|b{x
��{jFc���V�͏��Y9��V� �WB��T�1Ѥ�����v�#���rδ���_y���]�,��:�V��k�N����8�Fu�X�R��-[�nw?�c��JF�e�#����H���=�	C���S����:D�����4_6���/b�֨��hǻy��Y�"��+�_�X��io�^*St�*�]��X�m�'6�O����y+RF�=��4+�#�%?&0���kHn��|
�>G�,^�-�k�2������#g�&�%|eA	-�؅�ڼ�v��v�Z]�(g���YVʵ���߽B'"���%�3Rj� �q��j��^Z�Q^�p�M cE��l��Fu�?�ܗ����,E5T�~K���@�hws܊�`���A��D��o«t?�'�S,����:�]Ԗmp-qt���n�t9D�#^j�����#��ꆤ��HV�D�ū��CΗbvmX�A�7�fG�"�����CC�n����H��d�OGca�<��'�"EE�(K��Z��^�"�lb~��MХ��i�F�U�����§��eINX���D�ri�j������d�c�[ހ���&�����t����m���)��*k�����.�g{���uwaF\�k�/5��t��[�� �(:%6���`X���GeL�m{��Pj��S�:��7����e+y���$�A��)�/Y�CR�2D�
S���;T�Z��a+Δ�	֘G|�6ٰ �g�E	�\�g��{��:�?0iR2ҽ�w�u�}�=�C$�v59��4�qϹA\l/>���=>rK�M^-�0��ab	���,P��<��ҍ*v�B6��(ü�h2�"N���~��%��V�/m)��ϗ[�,?_�А+��9�PT��qE��������K �ʽ[=6 �ǂ�����{���g�����n�����Tۥ͕6���jm�Ð>�� [*H�d�SCӒ����ϊ��Жt܎�1aBڸ9���RD
,�l��J�(#�;S��ʵ-��}��-S�N��S�!���P����p�{g,�+!6Ŀ�����	�1anFA�زp �X*����FN��nQO���9��wx���c�b����%#��G&�i� 
���0KEx�x�W�$Џ��-wQ�ڕ���G{�}l������(�����\�����=��kB>�6����W��O[jt٢	�Ȯ�*1�mr��c��������C�CF�dp�
Ee��~����s����Y�<�?[P=a����c�lW�&=�	���x�!=���[�8�s4_�A&�����oDԀ�g4`d����C������<{.�f�O��#so��KL�.����l�
��Q����|��5hUX�_`8��V�(���������Ӑ
��^d�6�:�3:=�v��N�-Ce�q Qt$?{��U[��Q"26������3�k��u�'i��,�H_��r<E�W�qُǅÎoa:�97:$��	�>��HtU{�+���a�u�=9k�����h;ԛ`��E4�õ�ǽKccd��+شkN������������2-;�p��D>\��ں�Hq���'��lO� C��}�W��w���;�%HE���ƚD���[�0���	���j���[�h;�ki~�o�|��v�8͊쁆[wA����i)K^a7^�1v�q��� ��҇c9�[dU]J��B�!�|R+�@s�b�.�MgP,��0���}軥��n-~�C�bG@ߏ�FW�ilf�D�e�^3���g�XSe#����P}Q������6&��7"k��"<�(W�u��n�E��Y�^h�����K����z[
	�[1�Ř
�lRL{�g:^��d�i�anR,Gu���q�ib=f�#���@PZđ��eMa��P�n��A��� ��Q�Pf%�p��p09��O�d�h%Hl���rB��R�i,n� �PB�G�.Σ�X*J�����C4&Hq�'{덐|�k��� Ǣ�Vf�	�+.,�����oT�������G�J�-¦�D�A�(�^�U����	��%d���&��]�؊:�R��v6A�GTv�$�V�P��3��������ڒٷR3b:���<��Ė�&y'4����o7��ve`9<�7:��,Z�:��m�H�u�NrAޔ@;�P�up��7Sd��wQ$��6���Mw#������a�`'��-�nX�~����Y�-���x���@���(W�M'�ly]A��c�3��)r�qj4[�1��t���t}%�ׂt�M�[���R�gP�'2�ng��w=Ի���vL��������	 wԃ��5�^�ٝ<9є�U
d<�q �pzY����D?"T`���Zx��Ӥ��[]ԶP���	��#�C�U��ׄ����f���iK����7�CT�0%]�Bi���o?�M̀ /ݩ9 �aΪ]"֘���v�TV�����Ƅ)�-�=�ye,�|�%&MO�+�S��v� �Fo����b���9"��RϏ��=��7�g��z )o^�R`(k�r�$��uS6��g��ΐ7���#(%��}�B]��7b������u��8$��'�}<0��M>��C.�	#@�6	�s)�T<^�0x7I�rE]_N��&�E]��Z�
$�Z9�'���>jT�prk+<(Z�l�Ǩ0��SU�	��E���ˠ�PڤR	�c���0(��J� �M�|�9���o��
��,�����yb�diI�\�z��l���3��
|eŖ�2�pΔ,�/��lm_��5�vT�,���h!�V�~YU/­پ�����Ѝ��~�:R��խe��S��_5&Q>V@1CgK����A�?�~�PC�NγA���rjc"���T���k�Da/�Cjt��nw|0h�ަ�h��ů|s����癭N ����y�XT-��>X#'�(�\ �z~��.�%@�L������
�s�X߲	8*yzR��c���/��&�����^-���\j��,�k�MY�'�q�pɦ��}���MͳJ~�+ew����;Wֻu 	��pXnRGS�����8�d��x�Q(O���k� c�d�D���nЏ\i��pe�y���o�*}��D��b]T�]��ݵ��_랜~��c[�B���\$9(,���n��R�֓�t���q�r_�J1���Ѥ�~�r� �zi�,*�R����@�ںX\w�8zL���FJ<z1��?���
����C��2@��Wm���_2]h�
�EH
B��̔����L��Ä~�$��I��[�w'b�; :�MH\N9����s���D�C�j��	�͛$�-��`~`�L<F"K��[���.xŅ�H��6F�~��|)4�(D�<�J>�Эv�U7�����Z>�H�z��e]�@�m1�՜lT�%����G�?�j�;ƽnMs�WU��I��ıM���w"$! &�ql�������[�)�I��� ��d�ШXf+���z�%�N�Q�S�S0�:�6��Q1d�ť��k���<":����;���.��G:���|�O]*OA��������RW���M��g~g7��.i>sX��^٢eQ|�W���Ҿ�b]Wv=�T���[��*��S;�4!�V_��ԫ}=�^�L ��%���=���ֳ�O���s��ں�"A�*�c���2���y�ܠ�]�U��2��m�P��[Q\����9�2!Y��Ҹ�U�;Oz�����#	DKF�@.�KB�J�Ԋ����7�C�:9�X'�N��aKM����j�p��-��3�G;&��Wh !낵��U+��"�@�d@$����p<�W;�j��$�w`�D)0<��!K���C'"�n<��ly��L4���R��0W\"oh��ӑ�1ҿ�|�]1��C+�	��r�'��\{)B;��-��� 4�"05�D�W���M���k�N�96��6�Jg'َ��j�"���������`�KQ�a��N����$,U_��Hs�n��Ǚ��Hu=�^w�����s�5^F�߱:D��n:U�
�Ň��;K�n�>�W/�E~`���Z�t:�i�P���!a� \cU�y����Y��	6�	ETo�,�)1S��<���Iи�b�&PpU=��	���Y��x��ľ��㐛m�v��D��xV%`Z��Sqh��RIӝI[�κ(�K�:�J/��y�K��eJ�����8��εR�+��̎��F��q�R&�Y/4���.���?~�����W�<B�N�����f'���x�у�Zo�����Q��%b��%5���SL�f�0�+ܽ=�f�AlW_�°T:�P�W5;�jQ&߇-9">�&��%��J�b}Z
��P)F�����ƬZ���1j�}.������l��+�z$���e>�O��#ϛ�왼PaS�3Tɫ���F�a/잌ZyƧE;�����;'\ı�Uw�I�g?�JU�#�Gb�X� ���&��˻S���~\�x���{H�վ��E��.�Z�l��� �Jh0��%�H^�(������W���5}E�AQR;�H��̔�0�ּHk�������6�h��mj�����Bm}=E��&���A,��4�[㶎o���/����'W�t@��͔��E!�l;��������nal�"�ބ7���2A�F��5  >m��^�h.�:��8�Ȟ��z�`��H(���7>_���?҅�AUuϚk�!sl�?�d������y�'}��e��D��3t�.6�S��Og����X�<�K��û�D�#����+������_*�#o��E��K�8��W���E�$ZqZ��nb�V*:�p('����W|.^1�r��m�Q&'����}��PM�7_�p��{8k�[���K4�8�+?���{��t]�yg���5h}�ohV$�z�Ύ4O�n̲V�Ũ5�x�LZV7ļ8zo��*�D[�G��1~�GFX�G�b����Ҝ�֯����� Z3��],�N�6Y�ѕ�H5��W���I�����l
��p�'�#�F�Uo< rt�'��["��M	�w���U�C?ЮT%��qq�_�D��ʧ��v�M;�-h�F�l��{ ��uʉ=`2ꘒ@n�ύ��<��BT��>&��Ccq��Ϻ� I�'�T����p)�o4o]n?Q�3{8�J�����������R�[9��n�}�p���)oX�=���x�O��Yz�?�Ud�U�r�Yђ-1)|���1�ֺw���A�HܖFRހ����,�T�X�@��Y���k�3P�!'/�Y�"�?Ct�Xʭ���0\�>�Q̰��"q�
�/ʒ^j��c�d�)x6��e�n�O��+�a���w�+��kU�I Dng�y��PZ\;Sa}��nI,�j�ů�n�����F��ր)WU�KX�cM&���D�. ���(��KS�Ď�Q�{%�h�ѹT1 a4��O /��͝��S��d�����Hļt�����X'���eyc��Ãdh^��K=��r�Q*���T����b �H;�Srnk���\5�,� �|ٟ�z">�;�	�ު�@V#<~�i��@�X���/��{4�7�aV��l���m���4�Zإ� 0�������=X���0n2�=��d�E5���V�+�
�;�����P�?:1D���S�Ez�~ZT�s���u�!��(�q\��>�sq����E�rN.2�{\�\�!�8�P�T?��$��ߧ;�Xw�yj�e}�#�Uh ��F=�e羈n<�Y8�� �[V�Bm$��lG�kC.z%'�J?�g�\$Ѥ?n6є�:��󱉬����r��x'*��j����(���ެ���eF�0�!�9p�\'�j�<F���X�� zߙ�)��.4:�R`"iP�p[�c�-ZЮtOI�
ދ�~��E����/��I�}��ѧ��[�Fd���`�L����Y�#+_�p L��cw6�E���׼9�~�f9O�4Z�*�ɐm�H,;�ޑ�Y�!)�4�C�����saK�����Vg���6��I�WO���{7�NΞ?������Ov^X�j�K d#nSf#R�*jgLŌY�>&��B!����-��|:��	�=�MQ�Q"��~�0T�t�nl餴W���"^_�>��ۍ��������Q��j_v����d�97�
W�E����I�ݵ`	Q({]���A�(vV���b��e�I6�M] G�0��M��jb�D>Ŗ������n���C-�I��h=��^ZrOK�S�1�w�Lq$�Nl��Z�3��X
Nk��54��h����JG�����W�w�5����Lr�}�)@��8��櫹����K!�&��K�V�܋]�V4#�J�G��¢Њ���đ�qѭL4M=�&m[[B>t��.*龛�8�J�7)L5��~*5��Y`!%bs\�{�jK�?V����+��G���佨[�0��,ɟ���]Et3�������aε<�N�$���!$RX��Y�z���nKzj�&=לcK��ҢX��L�*L�`.�7��� �91�>Unq�=��t�[qZ�8�96;ƀv�T!�$~	_�穕IO��GH��T���jdӳ3�&�����6�B5'����T|9C�b���g$�ΐ1��Q��v�7���\K�
[^4W�!�[ t����. ��m�*��?][6V�Pt�к-�`�'��g�a�W�a���ULe)��g ZJZ����{�ct#�7�`Ox�C!"�
%�en��05=����G~^ԟ�'8�G%=�h:Œ�p����1j 4m�eb��2�Ȕu�i%Fi}g��]EoW��� v�a��*p�V��#���Y'vzD�EE��K��>Hl�Px�	2eZ��`�&H��Dݓ}~���#�&�E?�'3��%�����=��->��pPn�U<W�nA�,(k��TPb��˟(6C|	`���[�-拚!�����m��<�I)�)�sqݯ��	������5�_7��~�����@��EǎԤ���`��pJ-�hPY�a`
�V
.���j�#����	�y�3'�3�eq��T3�����~u�322�C�:U�3�g�R	��Ԛ����Q�>W������#ʮ�h5�VZ�f;�χ�#<�z>{��f?�#�C�D�J���H���E������|��x_�Q�f3b.Y�XӒ�خFWS	�C�������G�]+��C��T�>�r;46*gJ|fǎ'��A��7S��i�;4��^��.��6�%5FI�ՙH��i�X������'8�?R����(�g:v�؆��ʝ�i��J����ϊڤ�I�@�Z���!�s-u 7l�;�=�p^�:�H��(�3d�1a�?`�^��1�w�f��� �^�YĨ�C����ʕ�
ږ6dl��U�	>�����x/���Q����R����V�4r�[�>=x�@fا���&.߬�ǣ̍�7c�+�Xz��*.*�f��d{i\��v�rz>C9\�s,�EDeBh�P� ��J��ܸ{��"�o"��Rl_L��W�4�#�NG=�x|�����MOm�D�쇏����ɂ�ߝS���E"���x�Z������m�ͱ g�z?Z)���T��߂a�?��QZ�-�p�v������K��fL��ݢ@��g�& I�q�''ïG|�8��Qpc����o<K�ڎ�
8�Y��&�+����T���(`��k`$�{:T����}�D�#
�q#�����	�y�S��:v�!w{�e�}��4��e�BA
mwYZ�" ��.�*���^!�	�=^"�$~�*Z����fg�D���z�p�����[��Hl9�L��Ƀ&.}��MπNV$Ь~��咾s8k���RS:5
�}���KCUS;���Α�d�H�=�/`�[���ܡY��1a�{NR�n�@T�\���Tya�G{y[+����W]P	2���|�S�g4+b��-V�O'y�������_�ܝy��X ��M$�3��SW�yo�=��='�o�l�k	������q�)l�9;���
�7���i5��������F ��B!0rF{Ǯ�8�pv��z�w��O�VY�sOm �8�x��W�O��F‘����aҀ.w�C9�js�����4P� ����nRiҋ�/�8�\?>�#dnt��Z�n6m�@"�%���6��څ���^�Wu0�����C�����C
�D�G����E6ֽ�@�����cN��c �1L0)F�n�g�p_�V�v�Y�ƹ��C���#D#:Z�&�^�O�а4�b}^�ր�����tv��n��"\^�a��cUS��,���@(O0�]���Oh����;:���7�uxYAl�k�R��_`����1	Ҭ\���-�?�����G)@�?	��̃�n�#ֆ��_FB���i}�X���x���0|�'���x���!n��ѓ)N0Zj�h��ދ5F|#�Ś���s٬?��e���ұ���-��C�k�M��+�4,�NTR�C���/89��������j�� ���1��i�`����wW�����S-�Fn����aR�+-���vӚ�'��'�aȓd�8�|+�q:jt�?�%q�;>=辖b}�?�$�=��=�]ws�e�7 L���W.�@�c�7$�����#K��F��+D�Hο"�AG|`4{�+��b	�j���Kషȫ��]cOȇ��uĳG�<n�-�%�ؗq��/"�s}C�Tw/ �w0[�=��K�l�#�ԗ�נꜱʸ�XM��肙�pafu���:(�^c`��-Px0�|��>��N3#h��3�/a�V�W�}�PC��7:Dt��t1άĈ9�d�	оa#ox�?FP\0��G��ł���O�_C�s�2_�:]�������Z�DĒh������I,2!I��hF��?OnD}B�QX�k�+w��Q0�#!�4yb�l�nI���nV����MB�p���c%.��נ�E���J��{�b��	���P����-�!�+��	�(�X}|AD� ���z��Gp}���̾Ŋ� ��,"�O���Ql8Z��n�%.}�(24��շ��,��k���5[@��ǳ�j��x
&o ��n�_���I�КG/����t�ⅲU;"�m�R#<�Tl���ү0�5i((j��XN���Xz�=m_T1Ac�n����m6T�P�J'�0��A��&��ej
�pU���#�zS�Y��ۤ�zIѴ��x�#3���25�E�ÖKb�1��x@�j��z����]���g��4�M�ku�;��k���;��#��3�Vķ��`�Q��ViC�^Y�⼄ѧƒ�cJ���qe�;=�V��~t�H�����VzSd���O⟹n�O���}�
�-��~`ܵB�pMi'��|�ѣf�9�G��O��v�rhS��������+x��P�Y~A�\���\���-k�jv��T��'o������d��7/�~H�Z��۞$L
�}4�҂FvA�q��[�PL|�Yu�f|�XQ��x����;�P�")���)AC�� ����1�YUJЬ����mM=Q��s~��K�D^Z�4��l�x�P���L	�R�ll5d�
�l~D6~�KY�߭�=p��R�E_�9�%�����JJs2|MR^d��_����Ab����?J�=�
���ǳl�$�������hD�^��t���&)+�#&X�����n�n�ʕګ������&��7起�ҡ�[K4S{m������x_�S�̧ѥ�<GI��+x�o�ua�罱�HrBy&Q�Ѧ�L��ZHVuPPY�a���LH(r쎴<H8긫>WR��q�9�о��+����5���^�8��[��Pr�����H�ٻ�c��GYh��Q@|Һ/�0RIl"B@,�=�ux@��{�!�f��bM�KiA���{Pb3��z��[�:��/]7t\0L!D8��PA^\і�5/_��w�>z	cTg=��;�kU�ۉ���������_�"��<�4հ�Ds��WQ!"��Y��-�����_EJ���u��=m�"ލ��ڞdK9��&'qED���8�o,�5��h\���������N@
nI,�q��4�0�+޾���q�o�YZ2���;E]�����D7��7��]�� �JP��T@�|�ҧw*WT�F��,���_�3�f�����he���AI�y�O}�ۺ�(��B ����,���\Ɖ�`{<�X(�r��iqϚ��|�a�;TA���O�eM�]�[���fA�>�I�`k�>��F��#�6���PR}�R�W�܁{ݒR��.)L���������(��"�tr  u���;�5�q���[��e�.��=���O���JmI䀤�m�6-~`���5/M�OD�F�溟��[A������9΁�G0�;ɆGb�t��nWg���`�x�_~G�����Eb�w�(�'��L�2��b^V؋;��S�~��@f��k��ۋl�c�4/J;�����<s�m�=�`ᬧ����B���
��\jh&lS��H��ڙ	�>�b1fIR�؟��/��B�7��s��FFm�+���4�1�Q��
�@6ᯬ��:���k�Q�g9��A/+򿬛O�Hx~�o^>TR�Κ��}ɜE~���<�ފ[{ʽq�_şN�-S�����9�d$�q��䂖!��7��>6��ֱ�@��tx�R�g�.n��4�y S�vq� RMB=�BЬ{��
�샾E���
�3��[��1��R@�It�K{����H�.zB\b��p�o�`���O�y�Aq'@Ϳ�O�+6ҁ�N+��Ti�[7�I\�V��1I�0&?"��<3՗��Bl���O��K�~�N۱�7�����v�� ��ɑ,1cG�������g��s���\�%�6%��z��:-�,����`��3�H��>Pŵ�A�3��G��;?��mL<Y�`��K���z(�Not��R�w�{��;�|�{&p�8�(c+�������Y�6{c��a���gcG_>T˷����R#ĠO>��5�2�u,�U)/R*"��>�M�B4�#�W5��|r� �T=3��� y�Đ�ak'aJ
8�o��Y:�;6���q�=�&����d���6;:�k����)q!�t}��Nd��d�̞�ϻv8G��l���o�{8;�(;���p���3Y�GZg'1�.G�B�9��+�*�+! ��3]��ķ�j��h0۸�*�e�˒鉑iI�=���=(�sT�@3n�q���X�R�k{�+^�w��m�HҼ��"Z�f��ߎ�HO�:�V�/0ж�G�]�
�Ѿ��ٿ�:����<,�M�$�Jy��|��.n��`�������P��K�D�����&�
o6�"PĠMӤ�G�Lv^�5�-�$bo�%�4�h���"x�S�/�'GU�P�,������Z]�#�������B�(q�vkH�oң�qt���x���򠅳W�7>���"��Y�۪#-��@Yΐ$qZ����g<oJ�ݞӦ����pC�?!M�V��zQ��T�c<
9%����q�f��֖a�Rd�$�P�C!�	|�+�a��"�e"�%�g��ޤ�NЫ��4�}В�%`�"N�%�����|�PR�B��y�H~�>�4FoVJ���oZs\�Z_�?�Ύ����'��٬����
��@�\�����@�~�G�����a Q��4 �:r �?NA#kϥ4���~�Ӆa�,7�+����ĩ�ruG�]�������"&�o#��Ec[��(�Ǘ�]k��h�J��p�cH��8��ڗq�CZ�K-^�چ;�/Xw�$ ��{c혯�� ���,�F�ӎ��[(ĈJ�j���E�]\���f�_�I��:���E�@�y��6��-�Us%�����m[�h6w�3N��da�"��}*�g���s;9�J:�h�ە/vW�m�N�JGhx'\�sK���+���Jpر��!D���-WW�Y�pΛ���Z�>��J8e���^jr"�Θ��-��l���<�dAP?���[�j�̉�?����y�b���UgV���/�.J����l���:d=��xW�gҦ���n�PtL�&�9�
�6����~�1���:���0b4���X�!L�Q��p�G-,�^�]�j��0���w�N� -柤Sz�m3e�c���ؚ��E�F߄a�d;�2#;١D� (����&\-DA���U��3.��jB^����;�F�?���΅��FB�=���G�MF8�ь�xr�kB�3�S��ݼ'w�օa�dL�'�ӂ��������.�5��vF�&b�n/FM���s?��;Q�b4C�Ɉ�O.	^�R��3�O���n{1�����><#�ۜ�I�P [F�j6�tL"����q��%y��� V���0����X'��9��'����f+��p)
+硬�����#�C��\>����('��u��S5�,��qh��e��CF|�}�W�	
8'L�7iep�������+V�-��TwءJ���a�����=��避9i��ș���W{������8�]� u��^�-�@��՗�HrYSD��J��L5�YQ#���?�g��D��Jw���hf'8��;�9�<�����	i��V%*x:�	�WN��[iT����T�a�?sƃ�o�Ά#Q@m�Ǔ��>�� A&�ԗ�~��e^���e	�H���q�_�K�꠺t��y``ne����� ��d4 �"|~j�,���(P8����_���%��T����{�/;~���q�]�[D�%�ۡ�M�0Q*?uN���y!�����ߘ�� ���)�q�n-��y(G��7Ⱥ�Ks�u,�7&v_=Q������>1>l�<�W�
P���ԉk6=�lE��,�?�.<;��Rm"���ݯ�LU��0ԌZ�U��#v�Q{�����$�BG=h�����g�w�����7N��D�ڷ��]QJ��s��%CH��Ǻί���Ng����8[)��V`���ٱ�1ٛ�4s�)k���q���e��w`9e��2�{,��	1��=�_�S럷�əA��]k�-�	ϴ�vC
8i��$A�:���&���G�.�kJͷ=�R.BQ]�f!��G��&�y�!�v#`���	O��� C��ӾC���ۍ��5�`?�L5�I!C�k���;EҒC�� ��߉W��E����k"�*�h˱(�JHL%��n��ے�+F=�>�j0߈#eO x�fn�k�eR%�*�4��E1�3^�}��u7����{P&"�I8:�bK]�*{"l��k�F "�Yщ�5�aҔl�޿i�)�w�=��h���i��K�8�����=��au����q>�{ʂ�c��Whfފ��+�-��꿔�eP�c�O�Y�D6�y��^b��g�n!~�^��ΰ[O�B���,?�ӈ���u�s��F��_�E�dx	��_����E�j������h�+E�瞥��h�-�t�He++�n'y��K�'�2�v`�ݙ���	���枝
�_a��4��<�ٓ)���H�z��}*H��>�Hn;��9+i&e�3���H����E1�Ga�>@rK+��C�E�����WPb�X�aQ�H��#�9�
��Zs\RW��y��+����y@�7�:@�>���bA�pY���u:���a�r�<��~��k�,`�Sl�$�C�,r��:��t��y�a�Ng̛��m�����?@G\mEg����z�a���C:y�h�$x���f'�q/��dDŲM��g>��g�/+���
�_��\^�~_�D���i�ܬ����W�Wbk��5Q�jK��prNN}�x�P��_��r|�MO�O�
	�ձ��{ږ��6�����y��49��Q��TP����Z��׾��և�l_���wū����k�#_3��ɝ��$�Zv0���Q�����@�k&S��t_ť��;|��R�E�Q�R3f�9����S��9 Dq��nE{^d����c�Jر5�	�$��'`������[챉1YS[��W�r�_`Su�a�O�4 vI� �=E�Ƙ%��D���"7FMՉr��r18�C����_��B��3�'�`@O��-���c%�<4��[���]Hbx�w��㉀����'����|�y`d�$nM��B��AX'�:89��PX�Z||�T6`^@_����r$��Is
���!��$�1�Ds܀�{!�M�$�^0x��>cS,X���\#�'H���NpWV#F����fu`R<�ܸ�B��(�?���3���W�;O�C�E$q��)����*��q��D��`T�&K2[���A�X�;g��g YRu��X��kk)	A��3���"e�n�����Ѷ8��VWT��0�8ء'C-���M�
G�ߟ��>�L����l�VY��Q���sRF���\��5v�cg��7���Å��dH�xW� �)}Æcַ�����F�B�m)?�a;4w:��Ww���%j�-��8t�ElhU�H�W�B�H�],�����פ`	�!h@�dxJ��ڄ���3j�/�h�M�O���lY)ES3�Ƃ�v�i޿K��7�M����;83X�B��ΘѸ@yW����̾>I�6{ypVZ����.sP	��9N���؈���v5��<��V�D:�7���J�C>��ޗ������n�B�1T����RK����b�h~5FNDt�Dֹ�Z <��4>�gg�"�/���j�)|�z5Pe� ����]�g�D����oS��gV��A��pJ�*y�+���B��r]Q��
 �����!����	��n��z�?����b�ӱ�`�-�C����q�jƺ*TE>�oF��� _˄_�h���ޔsMn�b �%�xNw��;����`��N�$�No�1����K�c0l�	j�D\�iS���;"�vV�R��0��?;&�����fA��;�r='p_�%�Q�=��qG��7��z�=���@��$N�V���1R�Z$�]V��)���I��j���t\o�
#���
�p�=����<��?�y��t;!"�+d���|nNn���R�� �1�:�������,��G�̔j�bm{�e���>d��-.C@rhb�����n�(�t:zjv����Q��oc�z�k���"V0�Q��O��������$��"�g�6e��fo�BR(͚-[��/�(e�B�6�WՑy���v	�%o/�6�-e�EHD�6A2A��.~�Ey|wG�m0���������|܈�9>�A�V,����z���^g��m�P�%�+��s�X}�y'��:��hU�r�r���L��r���I�W<� m5E,��c([� �~
;�N���h�=�M[�r��|���$��%c̸�E$����]cdt{���Ȍ��eh�lLp��y���y�!�[&�P̈���;�Bpj_W�q�4}�<Ǌ�fފ��G���;�o���Fg�{9�R�EIU�j�a�k�����ң��v����:3�nqy"�k����}��-8>������˯��Y
E�C� C�+�h߫i	��+�y��3�L�(Ѭn4Nܝ�9N���ӫ�5V����W �_�ϽRmV��@���x@����;�/zƺ[)��<�b�]F6^0�u���4�ˉ
�w��5������jZ����y�_��}��Q%�'Ի��[�<�x��B0�{Ό�����AhJۡ��ζ�������NR��Sl��S���P�G�p�R�
�([��0찌u0�w�|r]{~��N�G������un�*\b@�����;Н@��n���@t�㓡_-4��Ɨ���z{��)<�a��-���鐶���B�뗘������ŕ�e�e��5\/.��j�V� �>�*��^�R�B����@V�����݄V���ZX�ߟ�l��������ӎ�5<w.��Y>�ked��Na�>�'�v<�����9$yW�w�0�T��tj8m��}R/�C�$kG��g�x� F=�?�=TOw�����Z��.�G�5�|�v�{�c�'��q<b���D >Y�hK�hb�2:nRX;N�����^��L�hs�b�SYʐ�({*�=Y?�{^���n�e[���Om>a�gݺN`t�"��u"gS����c�M�Xa�X}j Gp�U:<�/$�5��^N�=8�9|�e��P�m���χ��-t��X�x�=�Ug�|I|�,:���/��%M|�6U��UO�Hoه��ڥ��JM�S�;���p�)�R�����R^P<9b�lQ?B����M^M����Yk>�uP}�7r�����]�S���<L��%"��c��$&څ�Ӏ
��Bݽ.},S�ޕ����t+�ɠ�������v[KkQj/��h�|��O��K�� qo��B��_���/6�w!6xD�Wg?�Bk_-�ެ04ޙ�x��I�d/��u�⭈�dx��6�8�K���֕G�)}��]7�ke4��s �e<ľ}:���pVI��«�Nb�A�M��%|W�e~�-�@RRZ�*�-�q�%W(�I
k�3����ɿ@G�}��_6p��J��r�c?�_�M�+��޼�YB��&8��%.��|&f�6�_����j����kh��6k���n�Cwp6@܅���g�h��zr�5c"4n4+�.la3O��ד�K΂�<�r�Z�^73��/ɏ\�9�ߔ�k"ӎ�Ͳ��J�l�&xl�ۊ��#X&�݀�w�C�"_�f�Ն
��Ҕ'"�b����m��K)l�(s��"���`���>��=���,J��r��D��>��G����LI�C
�s#���@ڽX����$�**�弘�����������XB��?I�ź�YV��Q�L��g�2�_7�P׼Aq��{���+�WlF1q�i�ěy����x��@[���v�<WBB�ޛ֎?; �I���@b�>l%K|@V_;M�$��9|#�/U���<��|�k��L��s�Z t�95��F�i�{��2��|�uw{=���*�@u����Ev4�#Ee�m7@K���eiS��R,�e���V� �u�w�}Pkw˻v�갵q*��@�D�%<y�ٜ;�bڰ|���\�u��u˳���ȥ�b�u�1^Q+��<�ɌlQ�57�����S����Q��|1�+����<�~m�̓č9��ֆ7�6�ѓ^p��ږ�	��x��%�T�� �����ٛ	�v�	�f�P��	��#����^�2{��}�j`_.���?�v�#k��}=~�[�����j�G����T�ylM�kOJ0�ێ6��5�b����Xvi.P�rs	�L+��u�S�j1��:����Y�4x��O���?�ЦeK�}������RbԱݵF��y������>h��o�7cBǸAV�F����,�jm�h7�`��`t��x>�9�0s�++G�_�m��Nד�] ���C��S�zt�R��a��CJ-�CJ�Z��+�|���.Ag��/$}ҥ���V�p� ���<K
/b�M~�J���um�M�Y/�j~5N�^
�_N�%6M�O�w�	A�!����O�?9:3ÅV�&��@TD�p��l�5� шt$+����I ֔%��w5q[��p�S�RN��n��]R|�'!�a9L��M���M��(�b��_J�r�Xf��Q]��}H#���)!��k�)�1}���ݷa��679���Ճ{CRt���ΰ��\��/`��%
��U�D�^�
��"����s�(e�z�!��;��CG�w�W���Hs�����	��ys?2N:KY��%z	��^�L%,_�a�"I�}�l:H�󨠢�eNJ;s�2�d9U3=g�(��{���ȍ��s�Hӈi����4>�4���E���zc�O�#v�s�A���2�����w��l�2�%�����hV��` Y�����G*��s�o�[��fG/��T<��#�&Hu���X~ͧa�������&��?D�0ʫ�g�ƶ�+�� ����x�}�?I`w�L��E	R��AX_2Ȑy��y��۲��S����j}������s�[��I2;�P�T�K7Fŕ��W;.c_~��j��؁�h�4����oE��_��s�x��B��#ucŇC'��ׯW��t��"������
'k���'+ʘ'�sH����>��RN���o�\�(/cT��	*�V߀�qw�B	lwb�%���O��?�L�C�i�Y�Qa�wd�oQ@�#���� ��t�'���<l����x�j�v�)�O�@��"�E9�d�iQh����֭������{�$r�U1�'��<�,�~���a�&SY1 ��pC�?j�OE��=qژz��$�P��L�?��k��g�LS�
�k��6�����o�C|�^V��g&��=e|�h[ �4w�G0���E9���J
�x����>,%���*p�ER8���R�OVs)ࡵ�����>�+:��Ĉ��9 4�
���S5,�9$Ͻ��d���Gzs���h����B���E H�*��}����us2u�Uk��:�'(��4�%��Z�I{C���;̋�-�N<2w��������ר5�6|d��;�l�Qҟ���3}bOK͡��rhxİǗEŢ���%a��3�4��!|<�q��G���'G����';ԛ}%�$`R���itކzv��3ȭ�riq���+�AE{{5���K��Y� �q�Hu��}
�0
^��*�	i�ם������� ��%�'������fm�f9��!����ϰ��'����-r��v&�[���/nrh�c%���1�XT��V_C��R�V $K������=���)����u^#e�	��q8����n$	���b^�SVk���9�!J}Mփ����d�����%+!(k{�7�v��g���������㞳=i9�?�_�������]�$HrZ���.�u����3p���ե���X`G�Km_�=7U?c�s�3�kvdR��/�Y�
�$����$��y%�T�^(]dcs�S'ol˭��K7����d���£��QpM�y�5+���hF=�s?��s��6(6���ׇO�X�/.Qff���(n�r�Z��hf{y-��0z���K�Ȼ�^x�8�/8��M�*p$&B�ͮX:U�J��-�+>�np�W"��d�wQ,C�4Zit�gD���-i'?Vk���P���H�$鴓�2����$�4t�=�_{��\pU���Q�� LR�� �����:ݫ.�pi&���j�=���O��)	���A�6�3S٤�\�(��mu�"�j���'��D������s`�0����L�k'��pМ���G�
Gq�=>�/!�l,M���_o^�e�Ȏp��$��/&�k:ĥ��^��G�]��k6�C�ji|�m*C	�)��+�%A��?����kzL�p����=2HTDv�v�m�u���qwm(S?�o�'N�S�����2��E����U>@���<nX��8j���q�y޿90��x�+�*��vU�x�Ygv ��g�}�>����~%�o/���ɷnZ�v�)y��FOZ���w|]�?������e�TQ
�W�*���O=���b
(��_�_螣��wKx��>�*��.�����:�sN���7e�t�Y�T,�
�[�= ՜�d��HSQ�J`3O���y[��q��<(%��4��=���q�Y���3OڌWxU���m�ۙ��@�e
���X����<K/3����E��!��;E�N�RB,���� d�����ǘ�K�Wg�.�7���q�#:o2�0G���"V�M�e�}�S�2�x!�� }�����$q���w̝2^زk�\U�4�OY(��utV��!�ɬ�ݶ$���r��	�>��>oT0�����H[::�u|m6�����h�H����2@��*�� i[�XP�]���gy�>��`��U�Ez�6Oȏ���S�o|�)9J�CM�>C�W����ҹ2e�z�O�#��d��j�.i�A\ *���;L�hD�dB&���޽f�֐z�+N۠L���VZы���w� @�+�|s�?��3�Е{h�M�(�}uA�jB'?��O1B�G��E)Jة��L��&�����D�_]K�r�&�g.��\���u\�]�^OU
�?��	9� PG[U���2O��ULS]��sV�\����ίvfYG�KULS�[[���=�\/�1�75���"�����<�	���H�'p��9f�<,���(������/��s����!�����4����nR.��Z����	��Z�qM�>|*�:�����j�c�FK�����b�};�P�;)I�eYh�ڎ�0p&>k$����7�ɾk�:DAWw9�b]~}m�����|�ɉ@�D��8���<�d9�Q )��$��c.a��De�	�%GRW"o�\ �����w0�i�R����@�~�B'�+GG��bR��#ȜN��qd�KS�-�!�L_QD�W�D+��6 5���*`ì=�M�D����mڃcz�dW���$���gq���,=�����N�Efѣ�����-u
a�R�0n��n7�L����Z�1��z}r�i�m����K��·� ������BXac�.��H��8 w���¬G�`�T�4;w$�sc�r����z+����5:�J��;[N�[�Ø�?����T6��s	6m���v��s1�R
S�s;�tp��_#.�0���	����h�*���^����?ix��t"Г��[6�N���PH �zWIK���rt��jV�V�Z��Me���^�� 7���p)n�g�&hRZ/�"»�j���K~I��ål�dݛ���H�ƕ��9�����̰
�6F��1���{_vd�[p2Dj6��Z���>�=������a��%?��3�
�7׷�U�n[��HC}�*�%I������]v���g5�v-�?��8/�����o�����EL��Z�>9�r�=������S��D�p�ɹS&ݚ�r�l8�$�ժ�9�Mn_R4;vS���+��}�|n����{�N.l���PYDc��^�!��y�+��F3�-�k��_��kВQ4�-S	ߋ.����c?D'Ol*F�$6'�*u����[6����s�C���_�۝�&�xg�Uu
���SwK?���&;��#qy	e�QD�����)�Y\�ܙ��+��9at��:��|���7
�&d��Hr�^���9'��:ZOJE�y	�*ģ騟�u4�1C��d!�ʬt�I�p��PYuC˹�S8U���Q:��%�SXXl��(�|rmZb�1�	��f4�+�]���?+����/�Q�ig�rՆQ`~�hq`�=ڒ�]d�b7������h҉k��Τr'"z��P��c3�L@;}Q3�9rj��FY��qh!���zro�?s����,
�dY��8�`����!V�vC�������궩1  �"�� �v+�ܦI1�+ZR̨ra>��Od����W��XC�R��N���8����{������f�AC��?����}d�-�E��N^���q�5Q���>��vLR�%F��SI:Z� ��k����>,-��R�:��wi"E#��N�I�w&���l�W� )��s�"�S���:������U��G�:��I��7��Z�2�H�����~��8�@�
�	r�Ϥ����-�Asԥ��W�B&K&�%���w2҄	V�G��5 <��"Q�D���8���D/�ּSS�f���W�*Q��/\�M9~
�.D����l�C�6hM�9�L07�D��)��7JΝ�;�y���V5���bq5���ñ�דd�q�10`&����%e�!�6�0�B���S(t?vI'��j,��}JN��܀:��.]qci��F��S�:�跢�j�hT����x���?�i���򠦏�7�J�����3���6���lc�\H��Z5�	xO2�Mf@vM@��x � �U;�:-��lM'������,��J�z�"�rI�X����ŵ?<�J8q�z]s
Ҙ,_ȿ-�A�äc��z��Rmf�����uT�Ӟ[P!��>�P��lrB ���]��5�	J��*���i$M����@���h�VY�����V����'@~ VC&o_�b�e�J��Z� N{��:��E����jHP`R�dt��!,LV7	}��a8�(X,�1/6�A8������5oA����(�f<[<:�����t�"���?� MZ�&lw��"7����H$T�U�K8v��"�=24;�P!�;��3t�ŧH�B����><k=	�R gI��������Q�-������b�܃ ���;�A�|:�>y^Y��A�Y��v�2��8턮�3�G�mb}�G���R�f����<YI͵��s�����p����ZϹrz+���~v:;�
�	*6?�ϒ�2O|��g��c�.��#1��_w�C���򚅼dŞ�?l�zR7�4J�Z׍�fhѦ:�3@�"�V�����lJV��3O4i���i3���q�2�f��3Y�h���"�������i̰�����f�Q �����\!Yr ����4�Ǖ��^'���g��-�;'%��}�cN������Wz�ń�wEW�M�Y�u���[֛�t�
6��ƈ Y��u���ӗ�*�Ml�E~�\UV��ׂv��5��b�v>��l����r�6 ��w��R ;�-�[ƯM��{֯L��(Ϲ������Ӵ8q��H;;�N���N�0]�F�c�3��NU�j��H>���-%�~��&x �CSՍ�pK�|'��ֈ��UPjZ�S֩������� �D�W0�kZ<��ki��Μ��,�?q��5H�K_�`��)H9z�d��U���cM���k�G�x��na[�y��W��H�@e;��k��D�Ə8W��G��j9A�tMѣ�b+�L,uM�s���N�$�"S߷�D��N�C�X��Mpc0A#=doX\X�lt�Y|�%���7��?$`�Oݞ1C�yBg����;\�x�~��S�%[�Lm��}(��G`����biŃ�� ���l��ds�w����H]��yҳE6=լ�")[ש�6��46�e�X/����A�&,���ŧ��q�&���*�V�Bxˋ����㥤H�{�ٖ�A�|'$/�G����'~� ���K��ң�W�j(*�kݻ��Ć�͵��s��-��E�J�ma�R+^HS�t�}���z��lq�qI!��(�ր��F>�����7u�ȩi�&[灱�Vh�6�b9$�]�W�/#M�n�o���:��I�h��b�0F�u��daꬽz	'2.Ş{FԦ2|-�X�A%A��4Vx��h/~�Ъd.�b����5������~Z��=|�u����Bѐ�w��"U)l	'ʃ+6�t��VM�e�3�s��z�(��}�Gn*˥� ��W�I����O��dmG��'U��~�P�ī�/D�)�����%l�r�]�{e�^�4��㍚Rm��Χh�e�/�_fh�X�=�(��T�ZJD��r���k&XM��-��Z-���P�8^�ѯ�� �|iϓ�VfU\ tm!��jK��/�p�|��,��ўDү5���'��aQ;,�ts3�0��X�3��u��	/��r��˝W=�� �2,Lh
�ӣ7���K;}���������ʩ��# ӕi�;� "���ьA@�}ˉJ��Fƌ����q��=(���ХVk�$��"��WTL]TI2� �<01����R�yj'*S�~\�'��Ҥ4J��u	� ��.�#g|�-��f�j�P�C�#���?��F(���gE�GCZ�AgEHu�4�傒����W�������u��CCí�_|����@�c� k������t�Э����j�{��24G|~l�)�����ͫ�(�H�E����-����9�jo��ic�x����}�TK���)���1�s'�G�QR��Q��oܩ�����z�yq�������(�/{9�\,-<�;4B[��n�7*?�߻߳���Rq�����j&j�NܒV'�B ;�d�{��?F��L>�SH�yṦ�.�V�ES���p��g�K$1|�h�;���dG�o���|��AL��tW�g$��{O\7���l��Z����CA��3�,Xπz���^��&	�Wt3/��q��c,z�)Ro�f�~0go�_rmq���g��
����">���%W�>;������q�ҠP�d6e��K�-=ƟK����u�m��&���N���A��I�g�j,�UP}�$��_c�� ��1P`���ϋ������8���W�&faV%i����*�#_�kQ��^�~+��*(D�seolO�����D�k� ��/��H_r,��>�b�ׁ9���Q7K^ra�ClXX�\�Q`��ݴ~d�V�X�ȁ"���N�OVFd�z�]�%'93���b��J���;���P.c����Ɉ�$�ʳ�"�=Y8%6��&�+vQn�����<����zC�*��� �^m�����,����pTKL]�k��,�ަ�<^ݿ,`ӄ��%�Ts�w��mt(�k����K0�~������qV|� ���$/���;���1�]X��2���:?�X��>�E���C��}�:;5��	���������睁)T.�L�3c���Ku+��+�;����`5t�	mP�צ��͜SѠ4q`�Sm�n�E�C�_E�5��n���'.������6��&�p��O-�p��Z@��n=ۮ��}���z�S�������C݋=J���z'q��w��6I� ��ԗo毂}t���-�H�����!G�c{R�k�쎸�<`y{X�S�K�A�o$�|p|P}��pX�xQ�`�J�~t�ί�6|�x�ln7
�b���'����_��:y�������4M�Bk5���HJ<��$���V��H@�8�`g�M�`S��J���W�Ƀ	TZ��|���j�9˃R�`��+�خҙ��#���G�D,�o�y�sD��ʑMs`��+O(7-�$b6�VE���ѡ"qz7�#�P ���O�#���p�z׆���҄�u;vK�ۼ?-� ��d��H��&4�ծ����:��9�(�+�*��w�"~��D䠳�q_&p� �"��Ľ���ݙt��`fjp�6�l����c�����R��%�F�5���ep?7���!?��dn֬M�� �M��9��\�u҇C�t&m��1���d&X� �WR��I,}/+AWM`j�ƈ��h"���yks�]:ć[�3�\��vn��D�g�(;�/!J�\yr����WS !��b&��W�d߭�(M ������\^1 l#*<���#���)�OqҤ�ӣA�'����B�{Ȇ�>�hX�R(DtU)5Ĝ�X~Pb��2v|H�qw�(a(�p���@����h-P֦|���Y���!#���Ϗ�P�^a��%����7���s"aī�½��OI}Be�JЎ�t�����P�L�.*/l�������uF:�b�P'C-�K������6���]��\����o�`��ZQ�DGD7���3x.����􋙥�. 5Mۋ�4��B283�0��i�"�[��%�R�?c�T���f�k���Y�����	��|��!���4��K##��a���I��)�H0M��$��h�Yl���D
&�X����Uk���S�y;���`��k�!�PֆPI������p87��x��0IT,S���פ�G��b��I5��U�
�zW%X��C���#�_N�xvWT�Z8>$a�;	�nz�rO���-!>�S��ix�������F�9::��Ճ������o�-�--x,X1�k��J�G�*`w���^�����#e�n���+9ڽ�'�\r�p����Fu{\�Y�V�ώ�0sv�U{��͌����f(���N����p��H�����(RCZ:'��6։�f��]bL��G0����x�2T���&�(G�����4��n�}�J���h���}H(��i��9K�N>�yͦhsSX7_  C�mR}�8�]?0S}��� ��N��5K.��,lc�3lnMT۟}ּ�L�m�����k������f��
[�>�ʠ1���M�}c��CO�:���oI�<�/�'p��kUreaML��6��i�n��*|"48%��#4M��M1�.���9pyGM��W�h�o�8��e��0�r�E�)�U���s�"��7k �"w�^5�	S�$Kn}!��6�J1`eՔhO�cm�+�?S>}|KF�6��%s�	������b?n����m�yJD
��t(=��8�_U��XQ�C@u�	>��s?�S>�p�y8��
�
\�n"bx*8����E���J�=e�8�kZ�i �x wJ��n��,F��?��o��o�9Ȏu�m7�1��?�b��Q�Q���+EI�Г��3	�e=�bP)�B>���]ݒറ���D�0���!]��L�|?hkw�?|��p���3,^J}��X��<���y��F����ҁ �?��lF_QV�
 ~ͻw6i��Gr��uB��gX���E*����].�B_FҔb��*��S�����Om�	�] B�&�'��Z��v]��ƌ�t��=�QNsVg?�Ӈw��t��WKʊҦGgۭKp�/_C�ǥ�g$�7`�!�@Ƒ��Q=Ċ}��U�� y+��cA7��#.��OT�$�_�6�w���Y����2#�Ev1�,AT�O9H�#���l��K��T�ƍGeS�ఀ.��(�JJ��.�D4�ث��(� �2Eb.
�AC�Y���n6�*#�3Ikʢ����tǖ2�(e ^���t��vT�j�h_�׬ �Y�j��M�2�)ژ�^�7�-�=�(�H�S�0Z�ѕ��Y6?Ah�H��&0������p�����;M���\�p���X�~����f���{����#�qde�j�Q_�v*�{�#I�R��r_N�����E�]��n�O���G,�Qd*���D�U}0�����a���!��M Ls�W��������[b���O	�y��<E�]̠�h��Qz������֟�4Y�|(r���GS;ܯM�{���)
*�)�'�r��K��M9�������m��L��$��?��C��Q��B��=���zIÑ�d݂?`�Q����2��ƥ�c�����E�~�ъ|&��۴^������k!K�D�Ҙ���м��C\� ���T1�d{G��H�K��]��	2'|No3;$���4��=�֬��'�|rp>�/�����"s��%��9ڠ�P�#�3*=$�;�QC����P^�!�7����!��'�6�E,���]����|(�Wn���c3��Ѿ��e�|Vbp�N����-e�U�ʷ�k\���������~&�8�n	m]�%Z��(�'��������b܅�`6�/Ge��?ŵD��O.\P�h�q��^_n2h����)d�0.�A�U��v�ŗ8ƃ��ē}�j�{I��iy[h�;���Ѷ�N��1��'�i �(ӢYHHY���g�c�N(kNxS\#�Q���aw{Q�Q%�������.��b���o:[�b����^��ESJ�(�M�,8�;�����@�U� �k�����:f�q�Ҍ\�z�_(vs��\����+�"+馝��W3�V��P�K_d�5�iu��'K��?�U������,�RG����id�'�ZD��48�u�B7��1�BX~�k��D�׋=@[{�5}�9Q(���6�s;��';.���ʘޘ5��6ώ�������m�� ᷬ#��ոm�q�2�.��WЕ���8��oC�$�p喉t�s�(�U��/�e�&]J*���Ε���x5l�V�U��O�&#� mhn9w��~�u*G^��.��1*[ZW���?��$�sx�����
�A�yN�S��ض`;�D���R�yg �-�	%��G(�(�g��eJ"�,1���n�0R����'�����`��؊���4���D9d>�����ˍm*w�d��O'�C�ɚ�G��!K��cJ\����b��LBu�-��=��_ڥjk�٪_ٔ\s ��YA��,�څt/BH�p�|���!�5�.y�`6��M#Ru�bB�OY���	� )b������>�j��g�
@�%�s��?��\[�Cb��"����A����eG����,#�����!��cFI���i=8&�A��`�̞tH;�@w4��ϥU�}9^hbD8�C��V�!�E���ݡ��_����G��kz&������a�|�Dpb�ɰm��a3����s��d�l�2-*R�uu<Ǻ =ִ����v���s���"�W수(r��9���C��"�4,<�T.���M���RB���	G�/Z�Z�,��D��M��O���^`'v������Sa45�f��=j� Ewn����_I�슍]oݮ���U��S�ۀ0>nD����W�䁻5��4|���B��LEʦ��21,�]������k;�-��h�rG��u؆�
*D%�M�F*��� V���\322VL�w̔TO�;u��3"�w)=f�;1zo睤.`x�n3��&��ڂ�s<UJT/ %��^�k���e[��x�ys�,߭�}�=����!`%������UD
Pf'~�\�Gnm�~��"������ !h,���Pef�K����kD)��p�Y!�&$Cj���� ���A��9H��p�K]�����}v�p�ѱ���.<^�"��W��O�>�%��˰�" #c0OB�$�BFD�Z��N���(F�Q��۲��2÷c�c�i������#��u��ۭ`o�_����0 �/���  `k�������-���2���2뿛ǩ��/��x�Oa	h��k��Z�/n���}�M�~�}D��v�z�v�n��#�cz���=���OѮ)�œ�CKt�&�W�[�BX5��΃b�MU����Z<�Z���h���.F�J��w����[=�[u���2q�SN(�(Z7­�"#�G�K|���vw�7 2_�6�y�/ �?���B]m6R[�blv ������jD�N
��(�%v9��O�~�;ᯉ��Y5ʰ�����_�+�����#~���S{��R2�Q�m�F��/�$cQ�6yW�ʗ�^ӛL1*�ڙ���.�I��|�j�OB�?�-%Lz�Pc�%3ew�M^0S�v16��i�A-�v&�[AE�������&�ށ-Sߟ��O!���>���A��a�Vƃ��N�5��3=q�(GUM�Zb��K{�X��	 ��`x(��^Zy��>C�_��~�T��"��T,��~�T�`��g����L����ȋ�ZZu0njX�Dyi�s��%�s�A_����q<e��3�HMWrv|g|�$��>���ٲ1��B��u��<B���"��A����M�6F}��tu��A9�:��]+�j�2�9�"��u�E�����uV[��z�Ē���"�L�!��I^����[�q
-D������g@�#��Z>��R�o�^�|��۳ʒ�Q&^B�&�T\��G6����-ecz�[y��x�8�I���ss;�I�hD�P˖3�7q��}l����n`.S~��t�
��ş"�zv�CP�u�W_ǞJ#l�lv�/�Boh[�Sp��6w����0`w,9Y/�(N
�ߧ��9/��B��_?0�}�+�����Ld|�K����P�/�,��������E�A$N���<�U_Cf�O,�WԶ���[1�wb	f�w�C�����92 X�{-%}ܖ�z���x��4"��$�a��qo����s�B�Z�����`/C}�l#�+"��7��]V��
62��g��+��Л֭ԶF3���	\YK��hX���m��/�ړz';��MsY;*
މe��\�-�XJܕ�y��Y��Ӹ�z��tQ8�o��n��pM��u7���#��<a�̃-���j�hgr0���7��?��.:֧F5X'� �,���ܽ���q0v'���eG,�ޙ�@(��}$��#�<v� ��y<8]7�Yy�;<�Vi"$�~*wm���p�R���4Ŀ"^���'��X'b�,4Dl�M���$��"��pi�8S)7x�F�\\;�Z��#����O���B�P7����+����Zfd�(�����^����,(F�g���^k� xcL��\fâ������ '�d�L�;��V�ui�/4rnԛ��]�®��2���V�;�Ǆ�7�Ĉ �u��bEdx}����lS��5)֙�at7C=�Mfw�W��� (&�����%�E`o°\�U��鍲�nM�$x5I�C�0�r�>�:|#q,7��+<S�D�~���X����s���ͅ�Z���VR �
bXN��w�M���7D/f�[G�],�$̇S����>��\JMR>Kf)�5�Ә�4UO�&KOB.���� �~�s��U�0�juyi2���MȅpL�I��RI���3"�{��a'bS-���o�BV*E��<;^�7��۸����]^11�(�1]��Yxn
O.�Q��w8�Q�s�͋�����1�qE잠�f)��DC^��K��D�.���-%�!���l��Z�|ס={}7�8���#zI-,4��x�w_Ձ5֙�;��M��˳��$�ǎ�N�#��9(([Ι���z@��p'�W#�3���,�5����R�6��	W�`Cm�����
��;�;P<�C-�e��S��x��Ia�* �i;S�R U����`|9�Cj����5�F"��h%��?,[��0-t�&O�բ%A!8, zE����B�B���n���7(�J���Sv�q%��7�=����t�?4�n�{�������������8���5"A(X�ah�vy��_�A)<@�`����5�z�0Y;�IzP��g�V��f�/g65qvgE`Yl��9�fhV�,�����s�y���V��Z�gG�B�~�G�'��s}�颭s0χs֛�S�U�������СE1��H�M��R�ϫ�Yx ����S�YJ?�4L���zρ��jn�&:Zg�mh�;��*��RM[vP��5Of!�ʿ��\ŰM�-4<!��Ѝ#w���eﴔc�*�Ff*0n���f�8����`�Z��H>�EO�.��t��X��$R'�	�'zX߃�$(t�?�@�_�T�s����=>������&��)L#��gC�+���M���AQ$�m]�|:s1�$ݾQ�EXj]��we�P͑*c�A!(jS�LO��tƵL��g�b���-g`L~s>�;�$���'ګ|����C�)2�U����k*�{��'��KD����C��7�DR��wM85�`���P��(��s�Ctɠ�~�����	W�w~D��ΆFrT�>Ͻ���ϿYR]�ۊtB~�>�L�Yޢ-�M��\JA&f��|���'��Zo���a.���^/�+ޞ�@�Lt������2���k��,([D5/�;�%���0���]2��o;��4��D�9��d�gw��d+^�%}�%^���v�'�c���ky�'@K�tһ> �{%���*0�8�N�|lC����?�8q�X����F9CNC枛�3���}U�Z����>�Q��L�O�:�B�O!zݎÉ3+�{���#�bzs|b� �Fϫ� /~��I��q�j�M�?6��H�%?���c���A4c�Fc����D����������w���oVH-dw�5[�W�̤Zvl�� m#��)���9Բ�r9�DT�9���̊e8~��(��>��C�+��FK�1�n�7�(�T�}��*��ڏ7y���9e�3r�݂i>J Ν�����gW�5a������1�
�H�F����w�%� FT�9��X���b?��;�k��m�	�o?��@2G�li`�嵉��/�p�F,����E�n�}�*�?��XT��N��o��Q�A�;ɂj ƚ�/���JH�kZ���-��Dr(�v���[�Z��2דx�s���I3�l��� �64^J��I���x�#���	���Uˬ��� \���´v������O3�\�\&����m�v�qu v3�/��_Na�W&_��v� �tK��_m����Ml3v�'K��,b)W�{ ���J]LV�F�*Wd���Tᯗ�Yx�j�*Q|�UѺ+8
�(��r�e@/�aC�|f��>ƥ�t�	�W�E�S�G�������JDu���"�C_�Fh8K�_��`��)�n��j��{>�(q�u��#Q0��m�Y��Gg)c��YT>����J���i�W�ͤjm�.=R���,��*VS��yW���I�Pn���'�٤p�C0�H/''���c��֗6i�m��b��h�Ie��P��֦;Q�Lh�Ӆg'�I�`���2�;�UM��MŸ�pp9n���5HL�m���%��S��_?z����.�E�#�JH呮�f��g���Ι�zm=�z��`�Ki���?1�Ey9�|�꺖��L~�Sp�{.��!"ͯ�=�� �ʂ�p�d�6X2j��g�K�i�u�Jḱ9���&��{�K�cZ�g&�2eǤ�`�А3�L�W�6�4&se�*�Y��IW�Ƣx]w9�SfY]'t�����?����=�q�Q.e>����
��;��1ܶ![��r����!
@ɻGH�Gc�����zi9J6�Ĵ���ym�%��\#�)�t�P������
+ӍR��(�����{%|��.$��8��O����VM�"��P����h̃��ت8V���8����(C�Fͥ�X*0K�,<�?�Z10)E���Iq|I�>0��^�;Vt�)�t���EP�pi��$�[��A���~5�(��4��1�7�����~ܞ��p+J�B�*���]�Za�p�㋊Nȝ<y?ك����U��kwNH��sZ_�b��Ť��OP�>ɣ��&�e�Z&�,��=s}�zTک���q\y*a�0��s���-���q��.`� �H�Xj� �� ���M��:C8���>b���줟�{�����'u\���B%�-6�����g���"��@ܽ�͞�	��:��eF��xc����+��eq�Z��oϕ�ɢy��Y�0��F-$��x�W������Z:'
�uzh����'��R���}�ca9d��rUo�oY=�U��{�}x�.����� ����m�ja�巖p�g�\ߓl�m���1Me"a��d{��DB����<���g5�OR��Q�Ӈ���
�l�@Jǩ�J���J��b{�K�=��yT���0�v8�64�bo�эj���܅�ݹ��nD����o��c�S&�sl ��	Wk�_�`=Q�&E$Ro�l��>s7�U�,&8��!Z��~L���0g��ckU�y�ү��K5�4Ț��v���χ=�_ƌ�ٟ��̻���W��I���v�7W��4'�Y9�x�x7������^EN����<���Mrd�l� ��{òm��{w�C��Yˤ�z��bm(&
B_\QwS���v-��)�W\���)����i`tr�X���{*�ѫY�M�����"�m�������WG���A���YS��hOZ��_5*�x����b��2�Ű��+
�.[�=���"�ɞ�EN܁���}9�5j��Y|}4���KT
r,.	�]��1�P�	G�h�� b*�7i�����TL�9�����D�DJ���F)�C��ߗ	:� V~�_�Jx�����X(,�C1���eiH�}����x#���E:��x.���T�%�r����nu��(�[���Oo����o����@�+�b`~��1l�1��+ʴ �|:wЯ�������
ő s��ՆY)��a�7}�DzQ��F�Fe�,Jzl.�Ǥ��������P<91��u4H|�ϻ0�~�7Ki;T�o�t�*�i����6�p	�l�F�T�V4�y��Q�P��!����53A8K1r���>�yؠUn��b�J��nF(�0I��cI)���j�����*0y�5�,�����n{����BZ�e"��9L��2_�@��gE��(��r��]� c�?q���x�����) �z:
�?�恒��0g`�x"�PtMv��u(g�L[��4�2o��^@{�@"�
�[]9�Wj_��?��Ή>�yC���� �k32�~�S�7-�P���]��)̍��c�\I,����l���;��螱[0gb���k�B��>�ﮈ� ?�"s, L�z���Ҫ�����i,��tQG^�����x�z�N�ߤ@��Avtt֙���\g_E������&�� �(��3��3o�fIY~V�ѣ�{���K��B�b��J�QY��hu���V'����@z�%���p�r\��B�Ϻ�*�%M3��<�쒊��q5nBI
�p[��Y���t�づ�ɽ6XbP���0��bV����qP0�aa������=�f��Ӽp�^+5�m��#�k�!����+�;��5��E@�[V����ǖ��)�Y��/$��q\�G|��I�/QJ�N}ЉH�Q�`t(��{2^��z�7Ų���N�:?��T$9��Jܾ�=���b���5�x1ǇFEj�b�6r^�H�W�{?ו�G�/���Z'��GusK�d���ԇ��s�_��f��
}l,2|����vs�rW�ry�Y.u�OHC�r$R���w�	��k��$��_���0�8�E�.6EF<����:�wz�[�j.����d����̀,,tM�e�(�ל\��S��?�A�3�џ9A-OB�Tʖ�o|�sG�RpqW���� �h�~���ڂ=xm�b��Mw���5���R�S��3_3%(�\���)�l$����]�a3�*�`76��9�h�.h����rڸ��W��7RӋצ�#��R�������l�g�xS*D;�?�-�k�Ih/�uRL�[A����$�=�J�5ǐ�Y��5m��2P�q@57[�H�� �Fp��Ƒ89��}�qkO�k=m��d�ձ#��P�;$U�aE]l$b��?����6�A��$ڏe7��G��UH�����-^�B��j1z㢆+�� ��J��K�����PD>z-����h_�j�B�u6a�3�߀�5In�u ���ԃ�ZE5��Q��U�Z�XW���y��=���[Ӄ|�\���ג|>�`�K��F���۹�)�X��V�Mg�C` �#�]�A$�Tȑ�<���'!��%
A�Ю��޾N<vU�g�_�o���.��C�ƉƐ�6�y�M����t��F�C �^~s����S"��a꾢���H�[�:~�i6�/�Si�u�4EN>�\:�ZW�J���>[ޮ/+��:�Q6yK���
~������x&V-^,����p������Dÿ �SA�}ގ��\.떹@����*�H��*�GS�E�ҧ����߫�W9�&��Sn=݁�x����*s�O� �CwR#3�ZU����'����T�r�9�~��i`������^v�H������M�;�@�耭>�T�1s�b	�0�I�9��(O&�WV�D�rmhRۙ�r��P��D�� ��$âlf�-�B��v�K������&%R�w`s��.
^-�������Q ��N���lx�����I�7k���k?S�A�b_�pKT�VZ~�ąg���b���l:��m�뙅�&�zPP���8��'��"2\n�#�O�<�]�SR���ra$�q���lRd
�<(��%SJW��0������tIH8桐�ReZ����'����1%ÏZ`�'o�*"�?=U�~����nǵ���9WNw��G<e�r�<�w.++ʷ(���`d�*�l�[%~� �D@S:��ˢ�8��I�K_(XT8��;m���}��{������H�N��
3���ͫ��{ֺ�%�hn���3~N�IϢҀ����pʠ�z��ٯ�eV����%�~>�:��y]V�;#��d�'d��ж��(D����KWw2 v/�j��w��P����t�J^�>�LG��^Hdrƒ&����j�FVH'��'b44��T)Kw��"��/�
�k[��&Pg�&.3�ٕO���ZO�&�g#�L��z�خ)#C.@/�Έ�Ւ��@������ą}��;' ����(�S�I��k��j�B}]����ġ��g�%wTϩ��Ŗ��¸I]g�R̝�*����~��8��2�i�GI��]_g�m�t�o9��������ܔ��;f����@�m��N(��y�w�l��`.1!�l�~����_h�D��<�"��uB~��(<� ����,���u���H�!ύ��l6j�q�Zy�Po�Q���@�Z5V�z'�! �vo�KWν$���)��xè,������X�@IeY��CG���l��қ���V��K��+Zʚ�=����
�p��"�I��sB+����0. z�1���U	긓	�@��-HJU��N�4@$��y"�U�6�X�ܬ��;GCp������pظ��JS%����
�{t��ر;ٳ�� �>�kr�l��e�B����#W��3K�!�!=yzU�E�1d_t���f���?��ܔ]m�*�k���)��9���8��[�+*��f𔱡���o�U��e�Z�X}�9���/�!%L5�6�<�A�X��/���P� mwz r̆��2cK )a0hA��=_x��2���L��A� ��)ڽ�lf �⭳WF���ěW@Y+��y�/����Xxْ�k*C�y<�ɹ_F��n�%�ꙹ+���� m��c��s� x�#iz��dI�0�D`VI���b��;�e5�M��R�P�2p�Awӏ:܋P��i�/��������j���Q��O�䛡1����&B(�9)?�m�K��6Hq�>���*r���~tD�y����U��b�7R�e͟H'��v���BܸL6�?�h�����?�	�5����~i�Za�y�鲡c�%�3�ާ����XU���=:l�R2άD���;Pɼ*/1Sy��ی��Ze�"E���]p�Di%Z��:!�@GT"c� Ox���Rp8k�,�L �b��s!�xvTS�ˈ���;7������*�kVe�G1�<�g�F�?Z�0@zG�ԵIl��t%��R���l�r�R(]�,>X&M�=033�M���gQ�!1�:���C��t'z����n�U�o-��p������CWZ-
�o�&c�pơ�Ɲ�:4�� �q�$�a�8 Hiޱ��\��J�k�G;�C!�A©fp��&���Q���w:^I%��	a���RU�I�L�h��&=��VA���2Xm�����I��x��=� ^:�(䖝�8�ѭ��ۨ�.�O���k�]X�#��1�������ZA��;!�y�K��k�cw\����o���ܫ�R��p�g`��`���W�ű9q��uC��X?&I�1�46PH'Ƨ1A2�}�	�}��n^�q^�hȩ1	�@���j�.k�}�1-q贉�eWA�ɰ��@j�8��U�{������0[g�#A��P�N!ha>ĩ�&���Ӽ��h�! k5�a#�&q�����M���MD��_���Y��5�`��&	m��mN3����/I�.d��9������]L���<��o�P����4x,v�^�bQ��㸰�t�<�]�D�Cw�v�s(�����-�n�������Yc$����~��sUM���#R,�~�?{�5N@���_���=(#:VqKX;?�A�^�ԑg@A�߉
f��Q{A.�'B,��vE`Q�a��^`��Y-+$��%1�t��6���j�r����� �ܐ��8`����(,���G�����*��{��5Fk�YӎՠJP���M���B�x�s1BEw� �B���=�jej�KNf���ɌXխ��s�� ����<͋�I�O[q����Y�L�.5=�{@\�t)�$Q�lQ=��&i����5�RXXa=H��7:�D��K�����v����q�|�;9ϳ%1{�����@���O�R/��ET���U��>�����f�@%���#���QB�Cn����r��U�����)x�L�	�Ać��9�އ�
��p�g��KL����N��Q�����Y@ k���1��a�k�*ٍ^%k8������H����7I��k�"��q/�f\"��P#,U�{Crh�-�o�R�
�[C��,�SRĖ�A	�	g�8,/`�f���\�KHP� ���X�Y|�Nf�ly(�d�1�%s|a��)��{�,�����u9���6A{8,퍤���;�;�'�>���\�����3�nN�����D?�8�[�@�Ћ����>,+X�c������}�x��&'�r�X_��8K*��wmc���AF���X�0����`��R�P�S�W^⢨�7˙�5p��"�D��t�SX��75��:N��� ����n.|�LKA�v�5�:-TF^�5���B��~���q��e-�Gio����JW>�bĝ�4�Ò@	�͒^�(�����H��ȍ��r���_�� V��f�?�1&&jL˛���
���� ��Y�ڣ
�v������҅�#0]Ų�z����E{��qH����Sڡ*�4�ݷ��ZZ�W���B�m��}��)����B��)�z�̐]-�q�t���9CsCX�N yϵ�U*^�}й�Y��nv�9��ʻ><�sAV��Ez�(۝�	�1��sVl��=����	��!: �(���(bc��埓m��.�k�>�%nǽ{&�����dވ��'�"�{�-7U,��0�)kM���&�ۓ�(�ѕ�N�)Jd�A�[�~�X.峊��?�[������=gf૳*��*��&o������Ɩ|��І^)Dm^��!}Nۙ�]'!3����9kݚ�������v'YW�4?ihqY�c�34��������Ч�i�ͬ��;�ʊ���~�� U�V�_�W-��:ҡlu�I��3ԁ���w�$�����ߒy�#���	像��j��d��*ݳ�*��%�X�����G�³���׬��a"����� N9\|H���.|H�s�*
��H5���#���?�n�g����w�^��ҕ�{��9���
1cD4e��nEj��'G��d!��)�>��ײ��v(����p�>�5��� �}a�,r��Ķ0�,��	9X''��nu�Kw#	�Ƒ\{�G�坼'(ӮR���J�{��D��O�G׫��q7ۢ Hc���!#�>7�d�����&�8�L����hj_oʹAå�<��`�J�5���큶gu���pa}�`Z�{�Z���2+{���h�I�ǲ��Zq���t�
���9��sZ�����G:�N���,��S�y��k�H~V2"�aMl�f���,H��\�V�h!˯�j���=�f7ݒ��S���X=eʟ����e���,�E�Ѧ ��������
�UBO.`��m8s��T8�a�HS���r��tڨ�r^��'2��^A�F<��.G
��V'�,5�H�V@5�-�k�"ը�C"�,i#Qӳ�8�V�H'�~Y��[�{�8vF$k\��H� B���s�ƿ� �M6f�u���-��]/Z8ú\w
��ZP$7Y'ږr��w���eD��w�� ��?���~ԳWu��~�@���;�����ր� ����x����ŇQO���Y��}�>�M��[�N�H��W��V�.����~N����H�j$����U�����f%V!�2&n[�?g-��	d�$����Έ ���D:%wʥ&�5t����v�O��>��G�����ucB�����D��|e��&�Hhx�1��������H5 �V[_�>��
h7 !p��hSF1�ٵ���4�=��v2�<�����qB�0"�����mZ��$��I-|aJ�PX2q3`|B|]�f��扱��X��qs��ZD����A��J�w��y"u�z1��s�|k�C�f�2���N$��[uE��VO������ljW�o~����[�$j��Z��������Q�o1�M����]���-"N��4[���X{w�lm�� � �cK���#�[%�QZӋ{i?t:o�xg�+gD[l�O`o� ,Iڕܹ����ݡϭ�� �"R�=UG����e��{�ߊ��V!�x.��~���*}A��,z��-��]�����V�|C��=$?gQ�FP�[�������-���2��v�ָ�4YON���eItI`y�}M������>X�����?��
a���
.����A�Q+=��e�07�t�Y>!^>L���opb�(a� �x�rz�c�鋃��I��~Y�j4����{9Y���q�g.�i��K襽��Cǉ��M�Z�5��,����n��~�ݑ�4 ?�sc�-�eey0|%�I}�������Q�y�?.��J�s���3<�#8&�h�rRB���E�PH��<ar^u��Y ��ՈoJ�S4t�'��h��wO�@/d̞�����Y�E����#����<���R)��m4�*N��S�;��4<�Aƻ�mmW���njA{qe��"�x�{��r�����г�և`�Yu�Há(;^"_�]
4��h�jN��Z���4A}�Le��96�����<G�⺪Y��	�e���7�\�:jV�XA&~�y����+5�$E9�v��ʿ�F>t�5C{�S�j���K�<���)2G�,9��싪{d�-X��s)�/��svA�5�W	�����3�-oE^Kq@!���!o1�/�_~�@S��K��
�Kh91%,Q�/��~�֍d���������
CA��JlX����WT��&�7aUXZ�~��kM�Rʨk�����t��|8�M��k���� ���c*� %���'4�$g�1E��ܹ_<�U6��\ã�|H�T��O��[�l�\�=ʜ,HO��)c��{IP@ ����B���0%Y.h?��&���RJuY���#�v$��Z�u;{�,��$������({�LH&"��nb	S�A�-5+^5�]�܍>]�������<��unTK�>�iޛ���w��M?�}��2�\���(���5�%5=܏�b/M0��{d�>�N7�P 0�����)���D�X}�@�B��6t�Zf�/�t�o��ZU��o��o�uF�M�\r���xԉ�ӝ=w}E�+70��ߝ��(�?��P���M�%ѡ��o�,R�J&�c(Z�����=0��7B,G%�sVׇ,=�Ei!�fVb��4�V�񪝘�9jlr	a�l�>�:]7r���$9�`����Hô�5��W�y�@��^���S���a۫kY���u��8��pZc�ҝ��ղ��Q��EP/�;[�{:��B�̂��"��2A�pp�.����"�i~G���{�Rf<BT�!�vF=����-�#��H�'p����w��-���ye>1��r�-��GO�����mt�ӄ�Qu#ߵ�1^��)�zw 4�\�y}��;����������LN�f�-5�X
n��1�q��ޡ�n40�?ŗ�X�;�9�(��Q������V�%;��b���'�FC��q?/#�qʲ�� h�<jڈ��N�y����e����եnt2ω'����|��\D���+�t0j�~�u�-�w���'��x5����K�J�`�A}+�Ϻg���U��oԝ�㑂����]�	瘆̷��d��e��pg��n�����U�T_���b��W�$gNJ����ݫ���kk��P��<`z�zv
�*�4�䷌�Q���u�br��f-�+��������7��ɿ0"�bS[���"2�d� *��F�}D�S��,���6���B�n���Z�
3�X�s�ϤA��	��j.������?��ë����g��/�y��<k�e�Y@p{��(�D�A/,��A�b���1�xͮV[:+���M�[w�0޴]�8�#e����I�@G��vͬ_��U��:h�n>/F+�zb.� ��F�>R�e�}+��`�禾�����a�~�ow.i)*>%�&3���E�T,�.�
dt�|���tH}*G]6|O�he��D9���Y��d➭�އ��L5��c���y��ޙKd#��D���#5�S��4 ζg���VG�_W���ta���ؿ�"4�[����! 8�X�-�����B�����z��Z9���Ɏ��6��ڣ���F�����aS�t$�G��IVZu����_��Jx�x����Kb�ju5��I�@�w�=�;"�e�G���-�`P3��6狎.���� ��:�VZ��[����ȱ�0�:���{5��Zӣ^�_/�������B[�֍�n{�1{i?Fѣ��!I�s�1 �O�Ӂ��i{��0����75C`a/ �`��J�I.x�
��&3�Y�7�S;yP��L��)���: !�|]2��H�+	Q;�)��\�;^&��Q�f��+x����� �ֱi�&	�c�k�W'x#S�~ ��G[��P����؝��4��9���e��z�ę��`����_�]p,���kR`���*&cա+���z1���.��tɺ�$<������t6�gk�+��yb.kSa1�i�H��~�r�}k�ѱ	�� ���p��Z��RF5�6l�0�fM�d��V�TM�i�D����� c�.k|X�sB���EL�̦Oax�L���>F��ՙEȤ!6^@l ���BRpjbU6�k)���&��~�G">�Zl)���U$q��X߉��,v�b/�X�/�1:��>T;fy���E9V���k�,c��3�2^�c4ʚ���L�^ۑ�엄OmC��*����q3�Փn��n�/L$�#/������c타v�?���G��]����+ݬ�/��q�<=Y�7��O���|7�{�4����ؓ<~>� -�#�}!>(B4�x�� a}�q���T�����͂uM�VV�)������h�ok����i�ރ
&��e��c���`#��СX���}���Wh!3�9�[P�����&Fv:���Ie��ƛL�g��݃�g�B"6� �)Z.��=�"��
dQ����MB��x��U`0�m�"��ex?�x=��T��ɱ0]j���x��=܋6�9
��B����FƠ�|�"��O����y����D�I��Aj��c{�yɨ�!�iя����̅�1��hT}��M��ޫ��#����D�VqT��ۘ�̬SV7��s�ѤZ/C�)�
ƀ�u�$ZN`�O��H@��[GV��.��W˾C�z^�L۵�ˣ�]3����6,��(�	�V`w��f�LVu@��6��MG���n�Ղ� �Z��:)�ܝ�g�VQ��H`��w�F���Wd
��ن�7x�%y0g-D�� &~�����b�E��|- �W�B��c�����-K�q��A�f� ���������1"ni���v��{n}��:h���p�Z����n��݅�f�y|����f&�~��J�]���K9(`z�V���G\.�Q�ĕf�%�	�`z��9�>�5f��EzK�J�Y��h�5�uFܓV~ʳ�d/�1��C���,�k�ͮ��[��i�zZ+c<��w��K����|8��r=(3¾g}�3ե��1F"Ln�¨mڗ�CzE����e8g�7��<�ݕãñT��ޞ��[Y��=d#�p��*̃+��T����qFJ�/�$+M���Jj�0G�qM:v]�=�o˓}�xf�S;{�L<�6��f�f #���d�+z��$5�����1�@b��R"K%j��O��ܖX��M�i�j4�_��M������4�B�V��CV��'��ظ(�qŅ���,��**�O��$B�Mg�6���q�����\ݏ���z��Q|����@��n��S1epgy���j�IW�]u�T���'�@G���y}�j9%ȧ��c��DB<Q�$*������ޒ<��;l	�b�E�P�zrE�6z-<*D��k����3}��.z�u�X�*�yl�Y���NMX$Pg��g����E==�X����E(6�����'��4��U[�W����cĊ� 䦶��՝��Z�)�+�������Y�v����eƢ�5�L$�c�f�u'G�Vz��#%Sm˞�y�rb��L�����RSs^�Z���/�<F�7 F�p9���H8�nhB�*����h�Z�JgB��-O�0����X]���*샿B�L�3��%gA�c �v�ˌǢ�Ւ�4�)���$I%����g�J�#���@sV0m���09���Dt��2�"��ep͜�SɁxs;��O���ޫ�u�8n^yw}��$�/�.'��; ����eZ��IP���aC����P6j�=�2s���Uv7�]Y�blKq��:	��tI�8$����� �2��n<��n}�Շ�#�G}+|b�J!?�'6��.�Zbq(E��M�a�w5�-�+Y�J�A�UOU7C~�g�H�/�{P�42קH:��[�H�R"T��k&}���kK�)׷:�Q��Y~i��TxH�0��;VБ�/R���gz�_��dh���yv@�&��P��~�V�����n��~�i�ο�+��~��u�iĴ$�xD�.�������<�u�Im�n"l7{�{`��r n��&M��j���|W�-��F~M����
.U������h��ևg����W)�=�\��eV>1��
���O�ꭡ�(�d�[�9m'��5��J�Ӫ`�J� �:X���&עy\�qvuw�T"58��N2E�dP�a@wg9��X�� /[=�=)e�� ���
/@�_���sg���	P�#Aw�W�T7����'�g��@�Z}�9G�����c	'؂aWjτ�)Wj�6|F�_i?�a�]�P���R��1�z�v(G�r�q��+�J.�=�M�~BZ���h���Ǌv߽��.BVܻk!$����N��ws�CVh% �$J�D2u���r�VN EMa��'�߆��-�w�^�N�$�3�g߄O	�B}.%�K�����v,WP���l������F�A1���W����Ac�Z��[Tҭ��{�lk�U��:�6������b <Bz�Ӓ]��R��'�b午��0��&�h��/�n1E����_#W�h����wxt?��8r�92��^
9�~��`K��
�?�܎�b��w��9J����DJ���}q~�+�{���$���������&�&U9��b���v��2�Ϭ��vU��JEh�\����̴�@G�%�:P|��,��s����nUXic�fϤ��L��p��{NQ0QX6���ځ������#'إ���m0��V��1���:��CX��!�!��ڳw��b�rk�a�}��J/�	��	
��;<�%u@V�"v�U[��^ĥ�/'T6�R��^&����&�X����k�$����@x��s4��9h��?�iِ���L����"[O ,l"W�ZH��R�aXUw�5��`ڿ)V&�BZFŢ�őǵ;��G�t�ڴb@e��VǞ��}�t�ِy��"� <������vQt������_�.M�7���L���:��Ͻ���:�VFB�v����׾����0(�����6�S�^R�d��P�&����D	0:!`3���2(D֒k�p$f�1㟽8;����B$��Ҧ�Qm+��![�ܮ��esGf��@�k�����D�F7���9��Z�y�ó|�;�x��|�l�|���h��vv�|ZG�~�r�04\�&I�x�#9pB{�e�(�O0H*oTU�G��NWc��ty�R2ٸ��V�"����o���kĺ�S+31}�Z����`&�c��F�Ȍ� ��������{��=�X��bc�/����qbW��K�bw�R����j5�����x��=�� T��x�u����V��57�ƿ�*֩���\�VJ��:\cF�5��; `���1"솢��VY������of|A5�I;��f�I	��jN������i,�mj���+�t,��g�9o����H�x�!F�y�9�Me���NEq���+�p���v'?�`!��P�)lTQ�����V���y[r!����f�Ng�&v���D���qѠ>�ؿ�� xB��ث^��h7�^a���6�q�ޫgu�v/������3~���Ѽ^�9�ѧ�m��qY*�";���{�H϶�ͪ�ൗ�>֣Vv���kK�K4ͥ���:Y���20�w�K�(��#m@j�q�	�uDÄG�h
K,W��̰��g��i�fi���/G��r�g�k^:H�T����7z@�tURs�Ϋimz7�z(}C;G�d0,��]ԏ>�� �܋�ȡ@�e^�j�4�^���E��n��<lQ�0<�d���ĝM}nԞ���X\�!�`�O�f����"�_����❯Ϩ��q�(��L�`��o�`d��@�e�'+~�v��'���X�5m�v�;�� �n�-�]���0�A�1��ߟ��3�W��A�@�{T������C∳�*�����;o�|A7=dC��U���Z�N�nj6f�m	JV颎^�����w��<qD���)�F��g8�"@���	M�~�Q���c����� �ոہc�o��-��xj�M׵���I$�];.����\��+��m�����F��oM����=�1��L�,�]�GQ�9D�Zv%yS$��FMh�]��?@0"�D �ױD5|;ӗ�ø�[)�|egAdD,��Q�x��jnr�c���gb�0h��QSz��L&/�b�_olĖ8�	����a͞��mM4��<�	�:�=� .�Ԯ����A��@S�0]|�*��>��	A�v����O�'l2�yqc����J-���ߜ������p|~H�n���y��+Q�zͫ��}�*��� �U?���/\�S��J�}�W,��ر)-i'�����熜	�V����&�&���ۭ`���{sYp�3�8�����vM���A��zh�
x�'�E�*�c����"���c��E_��PB��tY�}��}I�����b,O�����i����e��T�'���z��{#?�h�� �n��c@�	xK����u��P��=�W�NL�
A��R��;ؘÖ����Mp��^��3[��:�	�uc���5��z�>A���x9r=��a��#h�6�Y#ϼ��FJ��
w�3F��ع��}�LE�&L�}��e1��[꾃�G�r��D�;�` ���s���1��|�ofe����D"N&��Y���[����@���S�����I���2.I��}~j#��đ)E�TL�ˢ����_��8�-ĒQBTL�t;6��~��	�x����%�R���ȩ�.H	�WA�L�-�'r��q���@��Pl�Ԓ�/�	�4l��[�Md��	��.��=�2[�����J��^uԯr���;��|F����	��$����Z��ʇi��b�>խ6���i���ւc���cΣ��%]X{i�'�M���/؛]� ��8ϯ9���Un�	/�:]��y�;=I�����7C-B�weg��aG�$=P����v��?�|�>eÎ=��W�J�̯������?(�N�;�,�$���v����͚m��K�-�ԔK��8�S��{ym�󗎌GL���te?��M܇��rc���%7�t���\
`�?;=�O����d����~�R;�C�rbQ�ti&�a�Z��`�:��%N�Sk�������9�M^Qwה;ߝ�;9>u�-h��Б��v�,��O��Ǒ�t�o��s��)����!ߟվk�3c���A�fW3�:ڲ���Z�j���cj:'�
R������sc�p�*��O�#�s�*ba�;�zJ�D��PG�mG"��[�r��E��!F�y�E���l� ����5" �w���I[;E��b�(=ǼժH����\qS琋�0i��2� +f��Ob�ԇo��KK����z'��/
�!�o������{�����y�Z3q���i_mk� eB?�2L� �<=�P� 4���fٔ�BɄ�{��Y5᝶��\�dD=ӱNҷ���#���ZՖt%�KW�`%�tf���f��Z$H���=*��p��� ��n�`��E�پw�n����x_0)�緵{أom�#Y!*2'�G���=y���Q��+�AkR}�Œ�Fl�ѐ=�k���&�=��`C�C�٣)�Ӊ;e�K��U�r	6�g݈L�����)�r?8Z�((H���S��(�Ι*�T,���rK¨�_��ԸJ�b`�:��p�x�_8����R/���=T���θ�=MZ�+.�i � ��(;O�9K��?e�5M+�����&~��{~w)�����̸�����E��Հu�}d���٪&�k��F�ޓ��T*�f�b��e>A{����]eCm6�G�9��^�vV����G�ڔ�;�4�����m�4�U�tH�F�%�J*-$�Է�(ZQr�u�兲i�:�{8������<ͩ�
`g8F����S�Xp��%�|�Q��J�>{�����>g�֫1B�F�UnH�"")G>�������I� ���8�V/nF(�L�_?�Ha�x8��n���n����3�<ċ7fm��2��+����B�H�o�����%O���Y��0%Z\�%71�	x���a �Mi���`�-��>a��4��Դ�ỨQ�0m�:)e�?xNx��_|[��#_���"� ���ȔT������N�'�ݓ_�-1'��(���\�kQFg\���t:�YQ,ӎ`@מR|�˂X�I�% ��g�o���u��\�ܰ����	��!]BQ�͓c?������~���R�W�q��w1"0n�PL��ü�Z��p���|YGƴ����z�u��D�����p��,�a���z7s"ﺬ��fWp��F ���o�L��V�~zD
OK����ot[���Z���~]�Q�M.C�#C���kU������b�ϑ��c�ON�2�Վ�ydZ^�;R8����9�	��]�t3y�.p���FX����o��a���I�g�����WqmC�nЄ�Z#����;r/B��5r����r�	�q�z��M2�v)���ŋ�]K9�`h̕�6���~@ܹ���y��n����6,��F<�B]Z�;�S��#�Y�e@@6������0��B>Y�y�u�ש�ާ�y���j�=�
(|2�~�s�kM�%�O�!�u-�@wf ����.�4S��b9 �S݅�}.�-y���kyN�A������VX��C�i��QW��/�׿�U6dc�Ε� ���h~�t��:��y`;�Z������ d��2w�P��R���K���!U��_�s�|EW�����-6����F�4nq,�S6�aL�аn��:��i� 륹��+Ȳ��6����/�vh��?ʫ��G�b	#kA\��!W�RI.A��s���HŤO�O�Q����~>��@����4B��K�|�=�:;�/�KO�a�?Z�'��[�0�űn]�����]=!����p+��?�*q��K�T��Pg3�T���0�wA�y��f��j�7˸�x$���u�cT��(��YU��ׇ��J�[-֞�cV����.�n
$���f(��ez�֭{�G@�ub�6�ӈ�|1�T�gР��.�f��D����J5��#�Pɞ�H�"�8h����Nv I��������н�~ � ���˓�����\�Gp،r�h��=�"a�0�t,���.��h&�D�^T�R@���6f(��Pe���@�~ϖ�#�xӓ�mwiJǆ�5�%�
���#8������#2�E�[�϶y�HA���c�|����jϋgБ���ܦw+�Ww�k;���}�\_=z�uc}�#�e�e��Eo*9�,Of�2�;�O�c )&�W���-ȝzy_2g��s5�#��b���h+��+=�,�"���w�������ւN0��Y��'�:;�gK��_��p��?`1����2*V�����Gn<D3qz��|gq��+F�|cW �E#?��p|��UT���tm���!U�m*��!�տ*�u�S�"����oNݺʓ~�7���Tj�̄u�R����Yw�?��';��J�YE@6=;z����W��Z�q�oZ)\��8��D,�a&��$!@6D��t��8p�F����� yl�����^���zH�"�KMN�7d�xnc�h��g|ƭ��g�q}9,�(�j�
���x�_�O��+�1M��N#WbΦ:rm�NU��$�c�&�{
�Haw�ED�Q꺡�����ՄzV������]q2a�d/H���x���n/��Ǆz1W�|?8�mG��w��_!#	榫�Q����)-��#@`��#�NL�K>:H 5��еX*�ꛐW�CS�:.���B�8#�>xZ��7$+P�(q���ķ-��@f���玘�8K�8��v^�9H��YJ]��â�U�'�.�@�T�7���	�J�fŎ,�9��p1���ũ�O����,4z:x�ߘIJ#\a�
\什�q~�u:1I�n#�ꐊ���ܺ���9�阳���T��<+��u;A�d,�up	�|*ـ�G� ߅-�i�Lsr�7��A+��j�ɒ���~�Lf�&���Z����cx%��R�����vF��8!�4މ�Ǜ�f��K'"@_	J6]�P�&@��7���B"M�����Y���CHR6�K���%��R�Y3�ȉ��j���H�g��Aq���v���y�@hN�Zn�
%p/�}HTǢX�H���Tƞ4i�j�ڮ��5�P�Ap�1F3�}�E�61~��6�I�z��,g׮�w���ϗ�ˇJǫr9�GX��H�f�e�i�<2⇲g@�#�]����qr걔�2)U�$�T�x�Ja�Rj�������S4��ma�M��e-�)�u��D
�{�5U�n>]�g��!҂�+�sH�'�������[1X�u��4��z�ȨES������vS��9����Ժ��R�RP6�*Q���T�\��٤�%���⒏��KFa=s�l�ۮ6��M ���R�;�I��~�F��4֒G��_2��#�?u$ �v��eq$���ZPWy�4�F�Ԟ��]Ȓ������0TE��!�W�+b��W�)q����s����3�x��R�3hJ}׶j�#9�DX�cM�{pS�7��q��{����v��s���1�U��c�&�/�_�������K��Y[W����'�$�&��q�/>��D�S.3.Ϋ�H�Cn1s)��y-�0$o��P�sA��tzU_\Ej���d����!OE�ݹ(M_����'IlE�}�u��x���H�cV% dG环*&�2]⮓�3�T5<��~�p}���,�/V��c��ޔ��uR4�ӯ��ti�%�6@k�5��Z�����:b75 �,ya豥u�LB�vנ���-�Ta����~��E8��7O�Sy�L�!e��e$��T�g���}+��ɔ��5{��؉P��r����E0� �׃�����OYn��ⵊI�g��!�P��l��-�\*N}O��=�Yu�ω��2S��4�l�� �
-+D�R�>��KM�i&�+����k|Sav^2D%r_D����$�iᵤx�'�~R��n��n�g���b�S0g�&�y�0�^t��cr��}�� ;z�lq}���ؑ���9�Z��~��8�]*fl
�3��n�FC��wQ�1m����M��������9��a��3Bm�����B����;~b}���N��-��2&0 "#�%�^FY�o�FU����S�ؽ���0�lR�N[~3I+�E3�.�0��s����b��=^\�%	�-^�g��WauCuʏT6Q�L�%�H�+����w�r�ɟ��o�u\ �g{������H59hp�?}{�R^G��ǘ��������SE�J��V� �U9��u�ˊ����M�E�@��U���z9E��|���'��3��Ad�a��x茛�0�"\j
Ht�wC	��~΀�̫��\�w�g��S0���<}-2�x#��MT�.(+�M�
5S�J3E��\Ɗ;�i��R��S�����N�n��	/���("�y��\dYĳN��L�V�3M��,�[*�}ɰ	���%���a��I+��������Ҹ����BY�L�\��ke4I)�'{�%5LV��z�����m�L��lU�\ڜsY)���ETL��c�~*-��x����o�'Dd��(g⅄��+�����J4��QP��q�B�P�p6*i�w�����c��~��d�{tFO��14�?&�,~� ��/N*��p�=E���R�،��r���~��u\�u��4�o�`�+�i�쏒�(����h�~��v/���S���P��cRW�0v�Kٍ��x�[Y��%�>�F�
��'4�s���u�L�(�[�@W���8A+�#Uj�m��W��ʣ=�&L����Fp(t�0e�Yr��S�x������Ϛw��2�z�̐����HD�r��C�l���.�{ib9�b�֡���[݊�
�J�������^q!��=Ps0��JM��J��S��eeb8C�s~�V�Q���>�
li�ږ�^T�r	��F�팆m��t����l�:�q�dl�sS~pC<�oA��������C�@�V�lS$���t��&�j�L���/�,~������S��"�	Yj�f"�� lW3����ң~�ɢ���J?H�Ls>em��{��s����)| ��H��o��"/��?�ci�%��d\*�2)o_�n��g�{.���|�������!A����8��� �E��4��`�{V���0]j�%�}�3%�I���!�Ň�������BƸ��ݰ:&���she����_�\��c�0�b�2
�PE���g���F�B��4��������6�l�����	��kH�]xCf>�X�� $}�uKva�ZE2�Q���5��~,(>O����$6	ܷ!L����U묉�=��8���rɍbc� �q��1
��'�C��n[�]W�����N��k�O�Զ�}Ć���p��%�C	{�I�g[�"���\�9ز3"7�q"��l�Q�a`�n�����Y�M�����,�ݚ���� "7 y�f}v��e�1/���]��J�Ar޲��V$b���вS��N���]h33�fw@�Q��s�W�v��J�Š:�B&n*'�����r&U�1}�f��۫���x!�X����'�l|�u��HT=ҏ�kW>�a'����n��D-�p�����彼hX?2N�H����g;�u�cV5�3��'^gJN���j( �z��j������N�3ЯY 0WO~�|����F��f��h���	%Sɒm�5�~��y�=�?�H��	�c�y�d��9=zē��u��4hǎ$�+]ȧ�|�Tgѿ0���T�������>�H������Y��"!�G�؜�	���Ct�Q�2�nL��Mݺ�f�d ���S����A��}h@��Ok�m��m�K�Y4@"�[;���!O�X�F19�i1C�� Aa�_w ������
��Zz�[5�$�*�uH`Єd�m���c�s-�H�y�t&���?�\�9U\�T��0D>���MF	#=�Hc�Q� �"���)�PwYX%��l(040���d��[�-0�� Pq���wsd���PKB:�;�ZU#@<�|���)�3m��+�2��S�����Ur8|�W݂o[Ɉe9hM��E��+��h��F��I\�5�3U��R�Z�
�O!���vH�,��Gٓ6Kg�JnS��~��!���K��n��%
Ĉ'�n���Nq�W��K?+��x��Ă
`�h�tl r�nװ�ЊB.i�6s�b
؜&6�L'�^�)#��ϰ9J���Uxk�(�/���1���^��s�S<�p�z�b�oʓ �p3����^�&�K�X$L�`P�&�E�Fɜ/>��.�!u����I]�t2�����vW����$չvU|����7�E������3} ��P��(y��AV�ϗ��W��fT�ζ}��]�!���y�I�� {�y/@�%|�����y�9��8����u]XBp,�*K
S-�����{�W�ư�YJ������!g��Va��?�f�;T|wk9a�^��"C�]9pk浘;y��MZD2Nf��2�����5ԷGE �P��Ob�d�D��L�A����;��33���i�H�k --�S'���]"�<[�
���l�y]vP��s� ���i���K@������a��)o6{��=�!��Pz��,F�0N��o4$M,�3,ַ����l��ա�;m��I�`����>�BQ����Ċc�w������h�_��W�DR�]T�(�M/��������-U����I���R�+0iM0�rfz��G)wo��g)��f��a��]>�4�4F 6HE=Lr�a�<�е�3 k��ܿe����|��N$*�`p��Rߦ�5����{#����S5�����o�,���.�f������O��_�Q�~�.�3}i����I�!�H��T��[2Df⨅aN�{���.e���ܱ2>�yŌ~Ŷ�I�M:~��XB9���-�>OW߼9��ۊ�h���>�KK?'��hs�� M;�"]�>�6�~ �������!�?�;��>%��#)�2�����\�+�C��z����+�zw=��>�i-�x���F ?O.�kFX�;���J���dh���c� �%�ۮ�pZ��� ��bX�óDm��a�~�l�D��ԯ?�2QՃ��#(�Z�>���f�<��i7�jXXZPU_aL���>ߌN|�Bqq���������C��D�W���"iš� ����>�W��ZY14��~���.Z�n;�v��T��U�O��jh�6h'��+ˈ�nL����`��3\����O��o�pf��pR-�?�Z��H�n �j4vj^}�(/Aj��#��V�>.p�=���d�����{m{��zp���0i�أY�(�1ݹ֑IU�b����Je6z���"��4k����6߿��֓�o���D����9����h�riЭ�׷3G7�R��d7��{!�*�i<��ո�2%��5
��V���M���D['�[�
��X�=��j�G��_]�i�8�j�Pc��&�t���	4�\ӟ�7j����jb��Յ�q~M�ٗ���b�y�����Q����d��4�|��y�V�3�[1�k-�\a�c����i�dT9J-)d~�8�A?1%��J�`��Em���!�}������[T��J�17�_).�&��K�@e�*:�. �ϭtkT  8�����
�Pp*N����:�K��J<�ֿ�c�;:�[9�<8�"�h�wJ ���1��R�0�nv0�x�����UMo �.�O�Kz�@T:m�9�c��*���c�flTAC�n��$ U��?E̘�ԅA�b\���\͉� ��[����t���ǶH�0g(�Gj��@����ڏ;�6��d�U���=���l�яyb�;' ��y�R/D�VW&~���N������� �y����B$y�"{=������wΛ�d� . 3���#�r�럨2�L��u�TB���}�f��-�?LE� y��
���/,�d��t#]Ig��~N�|:�U;�x.M����i��Z�BF��C�	��1�����}�4�ې~�� �7~�<�iH�t�Q �9c|#*А��[��g�Ď&����'?9X82'#{��<����ѱƵ��M�O��q�z_�UT�Ҟ͡��0W�f�S{����Z���zCa8�q��b�?��a
�[n4fx&�HZ	=�39��;�!f��� B��?���,��@��cM���"�/�}���x���
}�����юg��Jl	�M^�n�eqWe>���©z2��8�.X��N]�#��Z�P����ˮڏ�^:��`<F~T��}�� ��8� �d 8#rR:�{�0;���n/R	uJb��^�L�����h1KY��68�T �ʒxK�=���%�:�f���ƈ7���l%{I�ŖOc�J�>x8�^Q7�m����m:0��˼I6UtR��|A~��`Ly��mh�����J�ٷO!\��%��oI!�K���L���Y� ���:�#��R�P��-6�����d!]���f��C2��R����)����Q's��bl�[k��*r��.����op���3:@����7�g���.��|�*u*��B�'���o(m��>0�HS��^�b<" �ƣg�!W��Ƹ`�C���+���9���ڋ��l���7�m\pɂg���mm�lUS�Ll̘��G��r#��ՐV~�J3���Q�Q;�O�ʒ��iUC�����
:��&�;s�q��p��'�])>=��%C��Q�M���*��l~!��rJAp��f��Y�;�E���A�G\�L�l�D+,o��SN>��m�_�����e1���,h2�R}�@c=�*�y���{0��rH�\��K�� ��;�y�L\�x�+��j�`F.f��TDy�t������A��C�����JVǔ��Sve���]/�x7w��_5[�Ф�!BC�j(�F���WS��NT�ăJ�ʲ�{7h���%L&��?��� ��}B�eJ�K(N����6�+���lE���b��;vi�u6�3�T@Y������46�=:�u�+z�d1� ����.9��.�PA<E�,H(	�B9�y[���8G��-�x�Dp9�L�����wծW�u5�9cs� ����(|93��ۊ���o� ���m�K&:qj���h���bN�]
-�*'��O2E�4����:W���O���6�f"�Tp�}�%-!����3'���\95^�]��pm����(B�q�U
gz ��hM�V(2��G�f��se��=�w�(��b��Ol�C�ea��h�Amjl��M7�[��<�#eo��'�� ��	SVW�Y;�������P�,a�pU�̯�&
	�E���A8q������g��r1�x�Y�O	�2�ͭ�<�t�*0�G"L�d;��{���$@"0f�����j��k�v�����	Z����߯�p�	8Ú��[ҁ��|��eE� q�P��x�>����4?�42��8F��u�;.��񳓱T��dȲ�j���ycS����M�B�1C�Z�|�;y�h!��h���S���D�/�?Y\,�e���djn��ɟ�$n�mԱ8�U!����nW��n�$�P'�����7X rrn^���!�I@��Bwi���y
t9�EQ��F�M_L��fm�{)�T�DN.�ݩ�l(Gq��Bֱ�д�Y5��/��x���A�W/�4��-�i�o��bm���#a�Kc���n��;`f��,���q��w�l�؅m
����~�`WXА���֌���!�C�����S�������`3�g~��o�+�ae�fÌ�s�C��BP�f^�_ݫvT&h������#�M�L���6/�U����xL�����a�6j	v�ȫ��L�)��o�9�V-�gIz��%;�>}��KZ���'�H5R*�˽�z� ��L�h�.M����y����1�7��3�X�����+S�yf�$�^�·����bW˞�����`���F��x/�r���?n�HHĺA��W��FNe���ѽ���y��H��&�#�#b�3/�ֆ2�$�>`?�������I� �8 �%�*@]�g�@�e��T·_�R���
p�&��[-^�ܾV�K-NLeq�T��b�Ƈ1����+:�pɴO,T���wǑ� ]�N�\��i����]e�p����᫷)�>R���]����:>&i���#�R�{��s�Ea
����w�����q)���C2 ���C��&P,Շ`���O�"mE5x9%�Z3����ŉ�-��dV��M��R��<7r��g�~�YXz��ړ�2�YĽ�>`�|n�.:y#��hnʦ"��6�X�Qa�? ����>b(UZ�j�p�`F�P�\ J`0��f� $����b���9_��1�&S]��`���m�"� 9	Ni�)���Ђ�`�l��a8C�)�Rh!��rP����9�oBl�������F�'�s�]i%2��͆�1�=#[���.�A���:|��Wu���y�kc!|�)Vem!0�M*`<��7�s��d�h&�>��I��$�	���
`����2΁�����yy��WjhI� T4�6ٶ�ėEJ��hፍ(�ف�$�����3N��d���n*�N$���WBx�0O��������]������b=�̼�r���u��4���z������l3g����ev�2X������ˆ�Q�!��"�k���[Yl�Eu�#Q�l�?,!��u���?�0@��iB��A�)	Y����l1R��a���<\� �d���h����EЍ�7- ��)Y%�t�N�}���Ksn��
mҞ�ZaC��,�a�b1_q�	�e��3f��9�am�b��������$�3�����6�����g�zWpN�f���h��|��
n��(��T��pL��Mwt����ɔ�'�:��yv�sQQ@8!꬯�+'�pNPY�2�������[��)���K�������	�	�y�����'��\��,~BU�_ʻ����O&��El;�ߒ�+��@��,��@;��U8��d,���kw�u���[3�������ϧ(�D#}$��A,k���~�����vI�7����^��ahx��c��G�ui۔�����$�pU��Q��-opd��RL��҅����$�p�פL��JO���Q%�4����P���K���S@��8Qأ�CI�Ə�^�k�G#��'�P'0z�y,� s�=$�V!L��A�~[g�LR�w���{��������i�B���jF�A��ۦP�*�}��UWC�F�M��QS��	,t�P0�M�iC�@Q���2C�1%|m �U�fb����x�T���O��KRT��G'��$���IaRTw�)]�!�h\����)P7�,
���)�EX�\�H���`7��؅�}/d6�����V���D����=���F�D[.kK��a��jO(��{@(M�z�|N��Hq�K��^j��#Ͷ4���z,psG7SS�/��˘�D���%�u�Ll5���G�⍂��(m=�b�<�	Q*�.A����0��n.&��B���N� ꃨ
-՛��+4��`�k��?�0��K&�d���:�yKu"_��Ղ0ap�G[ǌ������i4~� }R�l@[�q�um��1�r�����3~�D9ɱ��$�GC	�6<�sHX=�����&S1�ֻ�
��Μt��ԡP�?*	{���[�,�a�_N�p��w��	}�H�1�����%
� � �{�|������	w���{�Z�oG�Q�Ep2���gJj�&�d����rKH��1�į�H��� ��o0���7��į�h�׷�)��� �u�k�ZM�;��n.C��n��:�Z��ZDMR�z�<v � �KV���0젓+w!��섗���H���HLW�ؘQCaX	��oz��]��1�{#��;�-�8'\Y�`����&�t�Qfw�gS���J�k�P̔�Kd��"s/|���"���s|h�Q�.����
�d�z�ꊡ����7a�%���<6/M����?�k�~j�$��R��B5�d}s%�(���`u��fB�^�gSe��SU����^ 6�;gcrgWA�9�:�V��;)Kk�+�b𸟗��ӯ��&��y ���V>�o��Ӡ�OY7�Ǩ����*�&��r�y�SQD?ѡ�
Ҕ%ƶ+�µ_+��x������;љ���o���,"��(W�1F����W��
��d�����A���|���0&��^ y	��jSH��
����t�"�LĘ���
��Ŧ�n���8ٜ�
�ؼ�E
`�N�ک�09{�Crt1��f/ �h�+�����қ;���T씵`��t�0����i>�<��A;\Z�U7E�2��4����P�$�)f��M^�h|p��I=�0��3�<(P��Ew��/\.N�¶��U��\���9�L|yU�P�4�O�|f:1 �ش� ����L�M΍�����7N�x/�y�l*�D|x@� ���GMh�%Nl{��K`d��Ӿ���	�VR�^�B���-o$z{?�y������ֻNq�.�L��-��&�MA�e}rNm�tK��y}�#������y'~���$�'���/��z�V��9PS�۾ł-��olw0&�u���!�q/���!Q�e����H�0�S^� 1d���<Y�C�R�����Y��]��y�i�����ìD�����}O]�S�m�fkċi���b;Z��aVw��,8�ui?�	kDge�бH�mN��C���3Yem)	����C/������V��泥�{ �)�4��TV�l3�Q >֚I�*z]����i�M��T`L������2� �d��]˴8η�<������"15Q�wT&UN	�R�.�3Y��Ϸ�g�C�����gLE�N���e&}�g��;���r����	��}�w)�.`o�)��ۤ��v��1��ųUԛ\��Jv̒j�W��,1t�<����X2� cy��Wh�u�t}�7>R�(���[m��]�A'�l�y��r	
��R@��N,�����?��vpu$B�`
�x��`(��D4���4�
��O�o�B��~�-�?�[�h�4�����c�$��.�b��=�>�]m6o�{F�la`�����S��#�R�"���ы�	��*�λ伿2SٝU��[��o�́�`6�#�4�r��q>=����cJ�������Ӈ&�0 ��9��Q�z{o�:ѵ��Rb"QGz���U�)�
��z���A�/.k�J4O.�i!.�r�RWw� �R�V?�[�,�j�|{Ɉ��{���+w���惎�v=�t6����se?��9Z�K���y:v?j��zΌ6�f夲*&��HW�W�3}��p����������us���$b�ɵ��Xn�H���;O1�C�fb�b��#{���<�l,h>�Riµ'�L�᧹�׵p�v�t~��ؤ�Z���l��6�� |Җ����Þ���Yċ��!�F&~���S}7��P��vث2K�_�"��?�=nL?вH	h��sJ��{n�W9_���Co�ϠfTԙ�� IF�0�/}=! ��`�6cOφ"��G�L�޺�ߦ�f�p��[� �S'M2�Ldg'v � s0��- � 
@���tN�E�HۀZ��(��qoA�8���,�{��D�(�wwP�+�u�����K���+��nA����%�~K�evY���8;��i���
#v�,���VI~�����R�^�v��JL�!����ߒ��ߖ��޲����䀿ׯ���[1�������G���p����� �&�k3$�e;���XS�[��:N�{���@���m�1a��7\�$}<kTx�3��#e���ۛml�8h̶�����nXqd���3���&-��Q�c^�䀸��v�c�Ukq�Dp I?@9�z���,|, ��lb�C�JAe�ľ�M�7m�k�U���1�=-cf��&,'�M�V��#�Ĝ)6&�ٴ(��W\`�ۚn�>l���&��۩�n]9^�5_O��b_j���Y��#�/L�؎�ճ�D�� �	<Ճm��><]��Q�� "h*j�Jt�?S}R�]�i����̗A8���pKm(��R�EO�קS�-ϑ�Z�~
p\�����D��p��=��CN�ssL��K���%����H�|]������:C�<_t_5�E�>�[�-��@(��mF��L��+����F)d�MQ���ރ��6�b�]�?�r �F ݂UWir�=�*��Y�,�'�p��Ey|`�U>�Cc䜫�+�ٛ��sz����kİ�K,b7�����\�����5�}m^��/���> *��z�-��Xe��'9���Q��e�_���U6��w���r�T���]F��m�n��Y|G�V���f�+G���f֫�yfC}��'���,������s���73�>,N�S1N^|��ʊ�B�֪�^����o:6�n�)^C?1�gy��H�Z���˵F$��v�!�>,����j������fd2QR��Kʶ��H���#�`�8,�=�#�2,&�=����Q�X�b�<m-�ơ9�G�� S)�o�T�8_{�z������%�ANj����HoWP���őwV�Ǭy��V�5t�~I�Uл��b����Xle���f<�L��8��٧��c>N7z]P� FB�=�a��Gظ���<�ф��ǥ����:U�^0������#)s�tJ�ᣗ*H�6�vct�?���m-���%�Cξ�<� �U�^��Z��[m�]d�ý��E��+������M��F�W֡D4�(A}MS��j��(rM��u[�f	�S��ϰ�n�jr��o�(R���4��N�wi�vP6F�6m-4-s�'�ȥ>Rxdw;u�h-<�v��!T��en�	���d�d��A�&�6��������&&��au52��������!��B��-�V*ZFq�k�q�>�@[���9�Z��1�q���B-+u�/I��2KJEQ������[/���XJ᥷g���6�"m|V��К�RQ̫BƜ{*��J�Lq^A�s*4���[��e�4��)�>2B�f�G? q����|D�B�`�54�U�m��xi˜S=��I_���%�cL��,}��� `�C?h����p����_���Ӎ�L�!����w'�!��E�ΣZ�ϣ�q��n��A�6/v8�������]#�_9L/ �F���^5Ŝ�f;�Fq�y	"���}L����ؗ���@}nr{�џ+��Ļ�3�m(>!O�O�#e�a�P�EA���dۿ�IY��1�ʊ"�CEƛ�U$��T�5w�n�H���u���nէР0�>v�C:��e�󟥗D�f�gQs�������j�p��$ں]�{5�y5�FY��X��J�|�$߿�o.o.�Y�#ӔR�����n���0"$l(T��?�R>k��o����+��l�0�C1e(H�:�ys���ɸ�:51!�i�^�"Z�N�|J�����p��Z�BX���`���@֖_n�aHQ��$���ľ���otZ�j�����
KKY�EU3ƍ������}m"�v��H�xbV��ٴ�v��.��qR`�"j���Z]=ܐ��%�Ob�zn�`����9!mzZ�u'��_[
�ȸw��!m��1�L'���a~�����@�-׹�!)/�
�Q��q�3<�����p,�1�}����;�Ͼ�U��]T#�1f
k�G�"��ʂ|��N�s��.�.������Ĥ��U�R`�瞒G�j]*�����b�2��r����jk?�LK'�3v���j����\�#����mW�1�[i荋^ĀiS�{E��>�u��(�r˟-�-g�W%3�[L:Fo����:��L$g'9����UчCÖ��xz�+����^D��V�M��=��� .��/6�Bʧ�H�<C���m�ph�10z��男%Av��,�`w�!�:�^����؄I�pVv�yj�tvE9�`�Uؖ�[�����|r�W�+��)T;mjݚ�4�M�U���F��Bk/�D����Ö������R����I�#���f��_��3��@K|vr��X�VJ�^F;)�zW�u�䊨3�&�p�u4!^9��Jq��AO�8�)�����,c�t�������ל�T�}�������SW�a�X�g>��˂�t���N������Ŧ,�u�DL�v�AR��t2P?�����
���Zƻ�N���O������NC��b�Ӽ��F�>v�.u�6V� rP^�l���<".�x0e��g0�����峼	��Tw�^9%�l�CF>ȓܮ^�Kl�|�/����]q���W��\�8&�PT���EL�NtOg�ΔH���B�{���Z!W��!�tb-�\1�J�J��P�6�QϪ��)��ĵ�~p� �[>�l*47��;Mm�(�<��C�_�P�_l��/������V{
J9��k{J��~Y7!$:���}�,�d�>T�U�l��DdK�x�Ɛ�n�~+�OQ=�*�V��:��{��\�@\7�a�<��G&rkG�?�N��&{~3h�D��YD& �^-c�z��:>�����w쭉�������D�JT��r��
w ����w��-A5{����A�D�U��=���מ�<˅�G�u����:��I`��28�z��|�0i`lG��d�;�^R��V?[d�_yb��:�cU�e저��5�I��ږBn�Ky��3�����ǖ@m�2�� 4^��h�/�ؙJ_�����v\BՆP焧�c��n�͊��M�Q���������S+��B�t$�����-����Mx��\6vg+����z�����C!#oK'������KQ�`����UxG�~^{� 8'�aF���M�+�a̟�Լ#�]��o��٭]�vz;moZ�#K��;�ܙ�qũE����4�[�W"�ȑl���%OeAX�K���eRa	CSJ�Q#[2�{hu�Z�0���7Q�'���c?~\��iGs$�5xc�[-���i�P�Rc�ݦ�%!=�ׂ�C"`��6�Fw̓f���W���7��� ur�c�����UOa 
��=�ܥ-�9�(��ڭ��N-n��IYg��:��,�a/6��?��(X�[�ymY�oX,[��F��5�+��$$���N�l`�t{B(�;�������;۸�!���]���߬���#A�ƅf⫉xYQ��5�U=��J�u�,mձ+5n4l(�jg��R3%C���/Wg��	�/�K`
�K�-Ec��6W}�)�x�쥁J���d �����՞^�fj�gbLBl�u�W�p���ʶ�^n�T3+(e�"v�&0����^cV��U뮻�C����g'��RH���l�5$����l�l3��BJ���m	p]��Oq�"Q��:���n�3�(&G��sRw��[E�LqQ+�7"��$��'��>W�%��D�:�'$τdƀ�J��g��c�-�C�]��Ɣ�O���4l����E�ZS04����ߤ	�-�GX�jF��H�{��w� �웰^�r�`"X��=8 |��H����ʓXQ��gL��� �i��r�?��x�6���u���{k�xx3y<܍� C�g:�9��k�Vkw�1.�v���%�Ĺ����Z'��qAM+{�N�c����/ɉry�dt�&����z�ƞ�}:1v�O��|N!_��z�?��HD/4���Ꭽp����g��p��4�M+ܟ�W����l� a�<<L��SNڥ��Ig<��@��䡷��"��ڹhg8dKݽ8�	�+>��k����h���}�T�/IqG�`P����<���r1J�"\A�	���d�%+2	+�=t>���^|�����C�J>B�"7������h���"�荍{�+�ăa.����Q�Fî`����>[]�0ţ��M��	��	};��	܉��eGy��8I
<���|���c��,�7���}��q�p�r�˙vcEqc�>,�<V�{a�%�!���*��wP ���*�N�5%}%?�9C$HV���r٠>�f�-����#d�*B ���n��o��x(
U�����z�"��Ϋ8�gP|�,`g�|$�/3�U��M���3���O_���3?:��qjY�x�1��1�]i�ok��� ���M���Ut��b���_{e�U�,��OKt@AB��]M��s����󦽝ڐ��m�i����ǝ��qfҜ��a���Y��^0o��>qf�ĞX"h�P>^3"R���i���c�LϮ�P��ﰙȜ�EAj\��>�=��A�oY��C���d�1��U��7�ܩD�o�^���]W �+�G�Q|7��с��t!���ՃV�������6m�ln>[��Gj4�q?j��SM�j��i���F>�XV�[��diZH���ّ�����n�{���Y��[T�~�\�XL��xJD`X��8���l���_n�@5pR�Nz�v�p�GKMu�Q�q���F�Y�Y(�I����-��Ǳ7J`i�d�l��w�~�=m���= .7��b%D*�^dw��Ε�w�b��{i��w�m�-U&��- ��?c䙥6�O�n�ѝ�Ǎ�MO���z�����eo'�L�+�=�ʨw�ɣ́}�q���>y3kٛ���eǍ��=ė�� �[<�!�h6����y6�rRƣ��V9D��'|6� ���Fc��31��7�\�;ޚP�X�`J��1��D�ʎ��T|=�H��0>>��S�:��㯍��%�!��sy��K��H���ęk�Y��a<]���m�)�(��窃�NS�pl�M]���U��?�{����I���ۣ��4R[�9)U��S ��vƤ���:�>�P�����n_�gV��M�!d�A_�WGg���������G��1�y,2�?q�����""[�U^5DۘB��PHG<�'�$��]�����	�>�zo��Is�Aj�߮#0&B�f������+L�V�U��BԖ�H���Q�J)���˴�?�J�g?l)���d;�MS���f4U���3/�\A�C7����H;X�j��嬓I��8}�w�%T�è��z�pE4��������Ԫ�0B�p5��@T��8�J�4��F��oQ�췛��ۮ�lx:�!���R�1�&�>F��+b:�z�Y�B��A���Z8�)[�Z ���\b�qrfG�%3��}�wx�n �CKQ
?�i�/v�4���𝦨8ˌ- %;
�z{K�*���,Q���J��5VB|d �W%�?�ӹ;-��kk�G��X6�D���4�|�܂@3 �1eQ�g!\)Z���È�)�h����2��� ����	~Q�di���H)ܶ����J]�Zю�w�~�sr��+r�\F����I]t�d�g��3NLGk*����b~�=�>C�����L�.��Kd�6 �QQ�]�2G��D�OQ-�:��&Y��*�77=Ǚ���{!_��|�E�&�aBQ}ހ�+�1�V���C��3�!Q%Lpl��_�{�I�m'�6A�w1��@)*���8�n	�B�.��Y�5���l�}o�K��(���$�� �E�bԱ%b�J���� 0�������Ft�k��S�l�Ӊ�d�h��&_�m�{�4�/��(?oÁN<rx%۸"�Kв־�yˤ�l��;M�er�Ɇ��iF�w`&#����5��p|9�q�4�[�0��o 5�	��yO�'���Oj�h�_F9����}��ҩ�
n�>��~��Һuz�N�6�+�\�����s���'��Ŵ3�2c��\@��7��!R���C4��L�Y�Ȫ�^׼z��F�<8���٣qLy�����fk�݃��⛸V��_��;fS�J���|�Q&�7�V��e���~J,d&`�^e;n7�b�}�T���0x�9#� ��#�'S�JlW��BN�jk���p�`��.�y�yU����g�� �-W{n�<��?�K��i	�����ye<��l�s���J~	oQ�Óc|��O� ���9Z�磱���S��e8��E�8���IEˉ{Ռ-��ZL��hkn{+���ya�A�8yP2��ऩ0�}�}���!=Vl�mZ�Q[��������Z+����B�bh��p�;:�C�ڪ;�K�2&�f,�h=yb�p+&�u��7g\BЖ�k������l$x���b� �~a�o�r���1��R4���."���M�ϥenw��q���!
D�O��	֌�܄��[ Az����R1� }ؘ�P.h�4�#9�{��]���vC�eӨ����X2���!}��7�MH<�(�# �T�1A[bຢ�%���{9 �{��a�pa�+�ࡗ'����NYfESmy;��r�G�����iLz���6��\����-.�������R���3�xd�P�7�b=!�����n��'���`Lb�Ko�nʁ��Pe8{�#P��ͷq�j���R6���m������D�/Q_�ؖ�4�K����w�"М�?���W��١%�^W��
���r�Y�#7lk�L��1۝��"��S� �:u}��x ��&6��s��$��@-~�k�s�,q8#>fC~N�VD����2pL���-*öD��W�v�);�
5,���%j8���$��(ϣ����."q��F��A&]C�[��	�o���h�Z��-�宑��o�j���+W�T���Yg.྅��T�]�
�:jD�%[bm���q�Mά	Y�!����Z>i۫�I�B�ZuV(+-)���]��V#���8��cg�h�N
�$�>u�"�g��A*CT��ԱT�,�*.r�=�i� ɏ����C��"F���S/ibq�`���!z�BL��m���&%���G�f��KǇ[��V�~-,<Yު�O�d}�[�4�����$�9�Y
y&��!$�D�^��q�䐎�x��`r��Z�����@�F��#I�ەJ�����	�5&šVkn��--�VӶ����i��<��#N�)
V�ZII�8|�F���?|��@��jM(� Bd!�Vt��d5-�a�B�%Q�Ȕ�SU"����+��i*���##@#��Z'hnJ���+�2{����T�Nn�ǻ����r'������,��6����.����r��N��k¦��H��	�^w���R����;�������>����B��D�ߴ6�t��$Z�ut��I���%�g�T�$���:'\�`w�����y�����`�j��y+�Q��J�[J��zr�F�K��qHq����H��0�Bn��_����u=��S[�>Uu�X�g�����n\�e�6iY�����H<�ǡ*��8|TGC�����ET����%܂ �V�0�`�z�!���Q�0�s��]a�f}恓�U���:W�Dfk�`?%�EE�W�?�=�!3��z��0�e�H�����]��C�P|h��cJQ;|���j�N�w#r'��"��{I���#�e��"�}G�rI]�V��x~�l!N�?9�|�ל�7ݙ�����W�Z�ج'&�2dG�d���O�]iE�'��K�L�4vY��ܮ���V�3_~�^K�zM8ߴ�t��.����+56���"SRq����z��i�a�7��zq�l@!�n#/��t���2�_r"&ʪ͵dwL,X)��)WU�\��i��n-~"�.M��؋U��5�=��Eb銳���Ũ�'��`����D�m�"g�o/ʌ�9F����塸!׼��fXz�!5ĥ3ږ	�<�h�	mI?�)@ �����p���G�-�F�D�1aI�i�'�Z`�/�U��� @�E�K��X���,X7�MP{*�<}���v�D�e
 ��PxC���+���5���[���ՙ�����r����ID�!�L�s��X��$��ǪܺO;uu=�Q���_x��������c�yI��>�q�lA�����i����"��.c�~T�TPQE�Ú�)�jZ"@�(��coQ��O�{#4Y�a*���iq_��Y�^d�,��ԵbԜE��}6\G���?��
�i�*)���Pf��TRe�P$����ڕc����H�h�����i�5��򸜅(��FW�.aQ��(�p ����h���F�w\oחU������AU=|�z�^�mS�C��HG��@�q�&��.ҥ����Ǚ;�Jdm]G��v�������;�*�@{J��j&S%����h�t�w���`�!]LXƟ"�-���t8<��yR���#�x@P˷�b*w�2�=5�?3 8&�2�=zD��JP���C�袾����ñ�A 4CT9�����9����4���� �y4�O�1�VU/I��a��2�������@��o(��5Q�΂Ij�����O����|&�sF;׸
*?�)�X-��W�tq�!7��K��؅!���-��~@P���Q����ɝF���ÂWe�,ܯr���s-'Y�Y=�6FPB���&�_Z�>r�����8.�]�Tr�A'�I	��o7��^��)`W�]�'þ�+34~f�MƠ��N^�-��G뒌�)���"�-�� ��+;K{��^��c��W�α���EV�$=R����=�ٴ���OjB����r��.��E�2����Cr�j8�gRm3_wۄF����V��\al3��u��`��W/�8��X%�/"�����oe����~��y@Y��ݭU���+�2��)w���1��E���jm��JK*�^��OzYȨ]뿅��wʨ�VP��;�IN�������S󧶹-�+�2~N��ߡZ�
�`��.E}<�Q�~�&�d���j�U�wyn� ��Z���`�B�8jx5��q�林�.a�s�>H�Cn�7T�&�3<Ip+����jeT@:9"}$>��!aV��� ��F�N|zPW[3�܆���{��V�Α���&��Y�e�������o��ԅ�[4y]�/��V�ǃ]xnl��>P��j��Pnȩ����P�_���A�'�����\���X�;�Q�-(��f����@=�B��<�^�����V#�E�hn�t��E!���ŷ�'n��1t���F��/���n�vQ���.p�}�	��D Q��<hEDM�/n�ȳS��N_V�-���M�Wm�*5'�߬��[�9�\*�<R�wN�|~s��uN�<�&2����v1	 �(�2�$��B�@4B�й����*n�������׬���̔$�*f0m��0є�Mz�;.j1�Y�bj�@��e�\x��K[@��(<��0o�=8B��Hǚ#?��?N�����]��4��L�0 .��-dS��@ɗ���9�/4޸�HhV�T��l��  �6�4��j���6�u���y����Sl(���/�q5xR��� 	�Ĕ�Z6��y���5�/��e�b���|c�Hg�T��[�H[��Gi���W�f�,�S�_�eCҫ}4���I�q�bd'	��l	�<u�O���'JZ����C��\��A�|O����@�֧3���.�St"��Jb�݄'2<Y<�J��Fq	�I��m�%�ފ���-�L��-����Q-0�/5j��BX�k���BG���R���Ǌ�vň�� ��ް���洖��o �kX�C�� G��������2V�7<B�Օ?�^;��++��-� ��[o�N-/����֬"����W����]���#�^j����֟c��a��ٔj����p�q����tl�)i2���Х*�)�qЌK�#�$P�c��	9��}t�S0�+��C}t��d_2�;t"��i��H����Q}�J ��<IG�쇠~�����n�,7y�va��wVJ����,�qɦ8��i
F�����<6^����6��͕C�RbL�x��"�f�{�������2*�����`��.�9;`V!�u �i	u�nh�}�,�l(�%F���S$Ċgܒ,}%b�4x��$�qi;�w�0T�%NZd�ǳ�qd6O���M���_XJ!U�yr,�S뵲�Ŋ��Y{MX�26��pKZ�;iYN͢'�k�D��C`P�Pf-u��}1��.�l��tNYyf��ŏ�yfL�:�w�v�E����"	�8�4�e�YZ��ʫ}vtq�	�l�Ջ��]�b�[l  ��"�8	��f�n��RT՗������{��;=�m��*��pɴ���8���{<\��
r���p���l[j�X<ï�a�(ˊu�g��Q����-B��l���`��Q��  ���(#�W��w�6�S�;�6�l���T˞�-C��*�ۖP��`���X�$R� ߧ���S���^l�r��^4V/P��%��P���G��B��1�w�d�J�a��5�V�,�~�-<��7��'��s%c�A�n7�G�A�q��D��r�L2���ߪ���?7���&&�S"��NJ�Opp���07�����Z�U��-o$K�Pr����qc{	=��T~`��1� �c�V�[o �ԯh��X
��G㻗�K�Ƿ��^��m�r)K�|�T k���ȗ|lG@�i$7��1�Iy+F�);��܌<�n[��#�_�����ޥt(�nVT������°�(���uP좟,1DV#j�_R�R���$8>��k��ףD�8�ȾM�Zo�XE�%�~�R�Gr�:�>�x��6��vr�5l��h��;��Z�w�ԧkKw'1�"�ަ'\ �Q1�?��>'d+k@T�4(pl`�X�@{���~
L�C�*|_�3�nw?~a� ��qg[?��,n�aC5�\�SI��Ug���@�מ�OK��tG�vvlw�%$b��87*�1�|2B;
 ,Ǫ�6�T�6lZGe����\8W/FGh�+3����(	�s�7یD�Rg�2����������l)d���~��=�`q{bO��{�%���|T�v;t�:��n�%U�QhV@&�1�܌����H��M��`�w��gk��
G_���p^�DT{�3���[	��G�R����ͷX�"<
��<�_��I3�ӎ&N���ZN��qV��Fpo�Pp�B>�axQ7>m���0b	S����j�����V!�_{�V)��g/�9�Q}�d�GB'7D�#<�]	�K�+x�q���I5C�����g��n��u%�PIғ�xY���nz��H�D̙���\��Ê��T��|lf �:�)�J��d�����;��-�=�=J�`Y(:A?+є��iN�!�#�V��p��2ߋ+�!s{$c�b�}�p��nd��]=���B�&&������F�Vmr9�'F?� CD�gz�|8���q2�!�
w?w�8Xԅ&>}���g����M����Be{8o�u���t�:��F����Tv\	��s��W��Qx� ����܆-(��it��i%�ō%����o�Ϣ��xN
�/IB\9W)���c�b*P�w����vr��Y�p�(a�x��y
�B�o06���l)3A׵&�I��p��޺S�n'�T��/o�p��V��iZm���?�������S�?�{���*Ĝ�9�# �C��T��AFCʐ:'�;���o$�f�wP�\�}�l�i��a5L��-y��ʐ&�J����C??y��1�����7#v����A�#��J�b5�r���5*vɯR_�nc�+�L |���όϩfw��Bq��y!��~	/l[>=�SΩM�~�������.��j�B$g��s�lqoC��9�����	�Lr�J5QWJf�5$Y[j�&��]X����!�Q�;�O��Rh��@Ay�����-��Z������9�G��b�t9x���qm���7��(1;wr<P�t+W9}�-MWA�K$|m�<������I�����!y��� :�:�_�+o�Sd|n9��/�W9�iڸ�Ԟ���,�I�U�����)�:%Y>o":�c��살�N�i�l��U����;����'!-�8F��(����d��e]������� �J��1e^�uv���F;,X������ ��L�(���$>���dg�+���BW�)�l��A��M��?�E?��6ك�!k���Ceb�O����-�t����|������Bqr���T� �������%�g��x{�������3�C��h�1<85�ڭjp��6P���#�;�A�̴�a���*SXw!"�$S��t/�v�R�a�CN"�ǧ���\wpjP�A[3�S�E_�"VJM�rF=��HK�Ēg%��r���3��H<�a^0�˹����SP�p�¶���1Yg��PM�����T{�^�;���,t�~%~&��qM�S�K�(W��--3��Df�P��n
����^M��#7�R��^���$�B��5,�^�n��G�Ypb����ޅ���J1�����������K[��s�nZ�o*�:�fl�z�wER=����g�	��F��6S�P] {�{�%nf7}mؑi����*r&L��ţ�����_x�hA�M����HF�RZ���M]�.�̇ф%W�V5�a=���I���ԯWrs���g�d2����s���A��"��
��c��b�,z��9\E��rb|\��Q�ڜ��ϻ��-�|{�K���Όx9��m�[���t��i���D����M����}T�)Y�l��$��QBR���X�姁�M����¤��q.g����`Osh����t�����E�`�ϒ�`S�촂�iۗ-���P���]�����Z���A�Ot6���*���䡵l�
��^����&'#*5%Mf�Ʈq�͈�E���w���d���)`h�6���yW�vbb���n�3��<v��t��w @=��Mr��2VB����T�N�hb�����B�#>�R���+_}��1A���,&� s䔋�';Y�|�s�� �-��%�uD�Ƿ����ۧ��^��h�9�>��@�J鮠T~�`��ݜL��3,����,�����bB�t���B�I�͊*�~�����-�*���|����k�_ϕ����)��٬,��Zc_������v9���e�~5�� *�H�1'N���&#� ���z@�2�ފ�Jq]�)�����*Sݿ��TS^$��	_��=a��a�"�X<3Y��8�����5s�&di~#�x ����|vOd��ʢɺ��-Du��Xǒ��7�(qmA��ԝ�in���}Vsϫۚ�J.蝯���f�
samw(ĝ'D	�9�F�~�YpMc>�Av(<,�R�y��ɾZr�h�H�a����&Y�)_�f�W�T��Z�M�6��M���v���|��`��C:���MG�F�wF�`�BW@7~����S�D����[���@�����t��ƈ�-
@��v�+1�ט�Op�b[U����(�=�R�ܾ�hY�����q�Sa2qY�H�c���h��ކ	�e/�h�c�hZfu�������K��J%ǂ��Z:��р�&AY	Vv��T4�[C�L�W��)&��f|���fY4c�5�W!�n^֬l�ҭ�U���Ɯ},���G{�O��+ u?MU���oڔ� ������!押4� ����W�k�U}�{�葋���N����a���t��X��c��2c�����Ό�PV���zS�̴�ݐ+Q��޼���<��'Dq�|=�y%���˒j���#��k�:< ���mL�2HvI;2�iPʮ/3��e�jd�>��c7�ʑg7�^ٓn�i<b�0�Q�"ߝ�nR���F���<�p@�h-�+�e��xP<�9Ũm���Xz:��Q��~ԥ���6��PI�h�k�0���~����π������>�G�
<��c�/v�Y�!�Ж`4�AÛy�r"d�ьׯ��(�����˨�����b�����m_g��8V���Cބ�p<H=����3���$b� �5N�j=�t�R������c9�:ʊ�~[�mы���-�3�?ײ��4\��7_߽�n�ƅ�W�%���僜D��A-�='�W2'�ףY��Z��m\��F��nl����k�3t���;�����%���i�L�	����z��C��h��V��)(�3�s��SF ���y���aJ~W�{���җ���5M�� o�ڣ�o`0�+9�ڪ����u�tl5\s[�U}V�������%H���S` x F�ƭt ��N�����Ӹ���o����C�������#��m�L��*�F�C�{z�N��mu�aη�\�@���U��N�|Swps�L�n�y����{�sHkS�(�N�]~4 t��4QR�c��9l��A�9��T1b'R�.�������l9؉�ʶ�FZ�[q�1�rs?RV�_uU��o�;�~S�z���a���7LV�E�7��q(�8][�=�HkѠ|�5qH����v�2ϖ��VlռN�����(�¾�>��^�b����<��O@��{���:��U�U��0�����k7Ӡ��QU2_�n�.��)t�����M�;���p �9�:�0�=��!G�L������NCQ��u=~�/H���&.VN��'�]���_�@��S �`0��9^��qm�E>=������8���.(ƻ���t���Z������е�q�qȲn���
�_|JK}L"�:��p���X�x3���Vo#�j��ܸ���_�Wγ-��T�KtR�rVkz�F��&�X�:��$�[Z�,WC:0S����^Ux�<u�)]�~�r���/v6^u�&0�*���1ϡ���,q�������'�Ω�t�c��]+'x��+�]��>?�jq
6ߡ��j)����Q��G�F�.��̆���������
�M{���F���a_�PH��'
�ʞ�8���gQ>��v��?�;,���"��R������^kI))��5o��N\�
���U~��ϻ���҄�d���!�FFA7�L٠Y�3=0�(s�c�9s�/�uw��*��������HqU}�&��<װ�	���TC;ofa�t�w��7A�������V���O���0�q���،����=ɔ��y�����w�kA��_i�~J�^��%a(|)�j:��\4e��G߫j��t+w}q[�x�]��s9�0ӌ��f��b��S���|E��$��Ykz�O�?ltM�{�N,�!�85F�Z馗f����vB���t�D�Q�s_�L��_�8�-�?Y��F������<�N����{)��ҘФL�b8��o��9��Α�'W�DrH�N�@U�u�0_�4HSx��O�L�Rݮ�����Z#�����m�<|�׃+�KE���G?�'M��,n۟BA@��t��n
���pq$�1,k�-y<Y�����񑜎`R�B���K� ���� A�!
�2(3ƀH�-���R���A�]!67~9�����Z�x4��7�lH���W�2�mު���_C���m,�3;��IR�R�܊ko��*�}q��&m%A�%Jz~�=�h8��O�u�s�}tfצݑ���V�Hh�ǖ���5��i���h��퇒��Ȟ���ϡJF��a{A	b��֞�b]F}���I`�Aȼ`���@�v��BS�߷2�v�j����h��E����/K}5��l���"�e-E�}ƒ.���B� ��p�6����S�T����3�R���4p����<Z��:jn.4�'Z\�(OL���	���S�����#a�&�׀�U���˲�TQ����vB[a&*�niWg><)yN�!�+')�O�X��o�_��v�>���7�����fJ���j� �/ӭJA.;r�
w0�*%IW)�:E�-,-�>귄j�»��P�ϧ��f�1ۖ�/7�R�Y���Q�?2�I�fv��1��z�Q'q��Ĺ�g##D5�J�0��U��K@H_�!���_��UO
���`K���1|�	���j�t��?l|3����-qk��T�:>�e�Yw�&~Ћ�V��8��č�oN��զN�
�ҳWHhy�/�Znk����5Yz%����4$3�aT�g��#�l��(��p�~�_Z��l��וBXW��b� i��}��ZOð��7���u
��+ϡ�-��W�n
��LD~VV�J���k��z;�F��
��]�LӲ�n_�{�u߃�Av��mg�=
�x��4�yE�B3����`�t+S��"?���Ne�k��X�
�ڬ��a�z��VF���&z!N�w���_~Z���HX�]T��[� !�E�#�OMƯW�&�l�%^ZW�[iAY�pM���S���P��k�*%E��s`$9%�4��-2����[�i���	��ʤN��g�@��1�Z���p�81��6%�X���&���~<Q���fřD+�cl��r�����E����w�E'	�V���AKF��݆{��+J�����	��I��v�����Q�o�*b��>�U^ܷ�=��p�E�X�W�ѷ�9�Z�n�i�G�΋
���
���M' ��U<����ŧrȸr�
[��ie��yK�P"$�Ǆf5�yW��yu��H�����UJ�F�9�E4����9S�w���0Hi����j�+.|:2�Va�B<�hs���D��Xk���^�t}�VQ0t��b�O�Sg���1K��:*4E��{l����#Oڅ��]?�Z�1��d�S;浔y2���c��>˛^zz�F(MH !jQ�� p��,K��D��'��[k���i5J��>:�f�K���D3c��������z�P.Ebך!7�}����6Ӆ���ط�(M��_U��j-n�(P	�G�oCl���F�rȔ�ݧ�,��-ހe�Ib�Ѳ��<��qu�63�ym�G/q����\��������uHbj�wo��Z�h0�oQL� d�$6/dEx�
�_hN^=��Lzϊ�b&,�	 g���y�	�����I��Ԁ�9���m�pS2�g+���½>q9�C��>x��Qk9���~T�m��W��m�d#����f�W����؁qʵn�a���e|v�+�!�#Ұ�c��n�G�O#DF����[2��N��B���z3�d��ٹ�a J�	��/��"���F.��p��P���818��䜫�(`>ϳ���v�Dc�cg��F��K�FJ�S{j�(8
`�ס��	k�q$v��C����;�z8=D6}?��F{�v��y}�<4�ϝ�i�
���[��"ĸ#����"�T�M�ջ�S��XW�~v#k�Z���Xݔ����l���1[E,Y4N��c����U@@�X�����GR�]���KI�1c��J'}u�U���l�ߤd�%T�F��9�g���.��H/�
�!�w�8��ɼ��Չ�b�	4I�{[.P]���J��i/h��n;�}2��� �#n�C���Uo��	�)�P�0��OUy[?�7_�H�?��V�(u���[�UH�����Y�}cyG�~t��׻o���Te(lp���	p]�_�-��o8�K��9�|��T�;o��ȟP|t_��ݍ&vF�ͺ¡�`]os=�!Ԣ�13eFk?~���-w�Y����P[�¼M}��F'I��k�[@��`���^.�y�0V��sM8��PY9?+�l�f��l0΢\��˴S��K��fM��S��,���tm91F9%L̰�ĄWb
 gk�����>6�%�߉`+qڝH��4��6 :��:�5���uR��/+s������l�P�D�A� c_ь��wM�Ezp�!m�,GD���oK+t_J�|�R�!��_��g�@ז�F��V�Kcf�oM+���cG{s�vG�(Qn�K��àƨv �&�8���+�h�/� ͵׏o^��eHa~��d��։F��!;+�v��-�ŧ�\,�6.���(JJ��qOTP#iK@v)�Slҭ��f�_Q�c��_ɬ��,�>̇K7�#Pv�;lH�V���m���_JFK��3�������W���n��P�g$�+�,�ܘL�Y�.'�{���a���CՂCc�YS�������re��2�����1�aFQ./mǃs��YQ:�c��m��p����E�� r�0�2�{�G��|��'F�)Ï�@7����-�7R˵b�����:�q4Pɖ,������x�hK*�-����Y��y�C���Zk��^�u,��k�(I6�/g
����Io���S��c0D����2V������F�����5�;)�̎prn��G�\m� Tӆ��l�Jd�I��l#��3�G^D��8Z�;�A���(Z�Jb%�'7�C� "4�d���X!sGLօj���1�F�!A�/g��:�oC�Gz�Z����h�����_�Jt��;7�����I�˙�b͸�S��G�N'�l��^��j8JA��\w�}�N���RD�հPWP O����N��<��_l� ǅ�k�v-o(��m��_��>�9W��e!�	�s&5�7*�r� *Zx"�Q#�<1�?�E���	Җ�z�3�]�G�;=P��r��0��l;{���_���d#�x^�"������<`3C꺤�S�	��`����N�H���"���.3��R3��6`�� ���SM��+�ٚ0�.��{�N�i����<^[�#�*��,Q�֩��	�}sv���x�6�~nFC�� ,�D��9�ϸu�a��-~l8�8�"���'$]����t�Cp;���6� ��3$Q[��G����s)H�y	�-��&4���夓z����2�A_��d�u�(d���2�JyXPЖƊ��zJ&���T�4G�M�>/��I�4�B�L_�謫�$������?x���ne��	��-�H@�-g�7]�x��~ ���%���g�c���_J��4�g����8�'	P��^��~��\S�|����*��͢�$6�LX(��?Z)/+�(T�~K���Z��S����e��
	�O�)�Hh���2���$c�q���&�InIC�U{n^_�.sİ�!��t��?��q`��5�Ц	&?�����ܛ��D?�0dc�|P;����m�����y�7�8�R ��F�mM,Ā��+lm��'H��6R�]���M�C��0���G	%���;��ZSg!��=�8�\*Eo�`�j�ghH|��a�G���9��S�ҞZ�?�N��ى���9>��(�6.m8Lv�ZS|8,hS"�u7͉�2o�Q�5EF�A;�?�� ��x%�Wd�k̅��w|���S	����������(�5\3
N�fN��K5��+��6����E�2[H��m{�Fm_�o4�V�Nk�nf��N�G��(r�u��F��r},�}L^�0v�W�� 1�ӱ�(衄(�$ap���2�FO������yZ�Imf�����xM��$�x_�rG%��xL��{�)j��.0m�g24g�&�z:HOe?�(�����PѬc�a�yU�)�0�<��� �R���Q��c�.�"�A���1�Jrᤏ��]\"Ϲ��*��-k	�.��h�&�V�|�no2��q��>��4��l��w���+ՑE`�!E�zxir*��B̪~����9(i3Ĳ���ذ`��p&2���>�ޚ3�Q�z
ݲ�e尓C�]ڊ=��`P�4,[�ma	\bHؗ�ͫ|$h�����JoB��uS7�.%c4�S�o��pL��b�-���S;6�E\���q��izWi�rp1Z�L�&&�r����n���f1��/J$ۚQ;��B�G��ୋ�
���}�ԥ��F�n܌ңR��p�2�ȍ��6���cP7N��-����E)��9B�?E��U���ޠ:F?R^0���}�e�t��.'��a�%�Q\�;�W���ԅ�K�Vi�h���x�m҂�Ҳ��w��Y�t��~�נ�>(�P�0ξ�iI/2��n���
�ɂ
=�p��y�Y�*��{�w�b4w��CAF�hJ@�B�U2�Ub�nS��]/
$�����ѧ��"���)\aU�7zfeZ��J���L��6v�Cmp W�}�u3,�s����5є���{��4ll}od���@H+�
�����"��ǈa2o=�X��<}�!�]�� F��h}t*�@�"��o�aG0���B՘Au=�u*(n�H�2=T���BE������<\*w�n��C?:��'u#N��1��dr�aH��W��=٨K�sp�n�Zd��zօ���r�EBw,tR�λ��dzӚ� �Ũ��F�t㘔�������V�pr5��ݔ�)R ?v��D}C͐�#,� �\���K�ߣh��T�b�A�.l�OD+��I璑�+~y�����S�$�m��W�� ���)z1}���Lm�b�:k��P{h]�V�卿b�Κж�nR�}X����xM�2��{�W��K�}�7қK�M�0���1+.o�
S�X�RTwSh����bXl�!e�~n���$�<���j,�3�o���/6��m�c�Z_!�l��q|\�д��e�JA���TK�`x������l��;Ŋ �_X�9������+���W�4*�2�:^ǆ�u˯��Qiաz΂B�����ڤ��2�Lk�ޅ�\J��+vb=�,��P��jn�� ��K[�#�FS�EV����.yE���>>���$��`t)I�]<t��x�iũ�J�̤�!��e!��	R[�t~� ��q1��B.�� �W�1T.�F�+�B���]G��
5Htn�ꌲ����������`(:e��]��?��7�W#���[��,Y��k��TÐ ���UF��z���j{�ۣ5rP�̍�W�$%�����ֳ�7&�x:��M�d~���[S�`g��1�ƥ:v^i����3G�V��ǔo�p�1� F�`��\�D�
QkSSK��n�|��8�<��L3`"���;k2�";x��0Lν�൫��L�T�ƌ�5�l�a>r,�q���7L�$`=4�W�Z��yT��bx���x�l�:P
�0�z��������Y�G؝M�"��/na+�	�Z��a1E%�,'�G����bş��=;��UX_�9*������`^CZ.wx�:j�c��pG�(��H��]����ʢ�%t�Vܢ��.�o�v���U��1a�㏿�P8`����J��Pӡ���I�堽?C��#�-պA����A:� �����eS�;�j*�I�f���J���UNբ��bqn�=>� ���~lD6��j�l�4;�DR.]Ul�$�P���r���`����i�G�f�U�Ӷ6q���M���K<�ɱ�I?��E�J�(�xߩi�[����2zήu0fo�l���R���c;*	"� ��ֺv�P�bB�P�Z����C�e�l���6��NS�(��Y���5a�5-�d�,���r��������_9�/���{���x,����V�"-�&�^�T��d��urtd%��
A�-xP����vϠb�:ܐ���@__�� ~�j��vI�H�M����ϫ�I�j�q2I��^kF���$Э����+�Ϝ3�\ԠՅ��Σu��dOkL1���"�0O�{�4�%# cC3S����IlZ傧�x��z����q���3C?`���c@�cs�c�4!��'��#����O�**1��9��a����iZ,!�Z�ғ��' VϩNR ��V��>�A���7��������g�G�4��n��{�;�TC{�ᕼWY,����@���Ȥą�R�1T�h��l�d\�)h���������Z�8t;n���r�`T��T<��'i��V-�}�ָ�4^��0�dQ�M�褩X]��P��K��S�3^x��_{d�����,ܓ��6Xt�Y������#	��-��S1�����?a=�Z�d d)�PB�����{��ӟ�1gR��P0Y��p]��zZM�+ �-	ѷϱ���"�ĩ��gھ&��]F�������h�~�#c�[��c�5�f�<'�E'�d$Z�6��NG��XW�OR�Ơ��,�rW��s��2"��l\n�Օ����e����!,�Lo�>d|_�k�6,8��6B����DAR�h�إ��/U� ���E�2~g%�2j����&��A	�,5S:�%Tb�S�����Q���x�f�����z����u��k������2�"i*���Bm������κ�_�K_�IY.խ�f%�Gwr����>�H�9G�����j:9���	u�^�UN��O"7UI�/@r;:�E��1��w��@ 	����pMl��Z�}sLI�W<ϓ��X�:��R�fY'�;F[{�%1� �Nb�(Q�̼vCToI�N�>�C����<� �4��x) �;ky����;,����)vG�)��=�U� ����\"D�}�������wI�!eH-�ubcvy��!���4n?����Z�f�˖ŁE�me§J/U~�	�m�;d��K����9X�Ie��%8ɠ��/6M�Y\��\a"�F�����p�\�3"�T")������y.�=���s�)�*,+X͕�1O����~�����X�X�گE5�-6��55w�=���FI�'^�<A�u_�;a-���SQx;�4�8M�#S��꒚��˹]t�j��BO�_�$�ma��"R��br�^���nՓIѧ���SwaK���f�=����	�kMt��c�jnV���CU	O7��';�v���͐UPi�4?���M�^�U�5�C5�`l[���?���9��*��N��|���@��GF[7����-:W�=����ٕ�Y�r����&����e��E�C�6�,���ZsÞ�i�S�ƥ���������D- � �#�Dm��0tY-�Ļҋo�2`U<�]Ph�AJ!�@���b������uYu�`�ww#t,�JR�:6���T�ٶ;_+R$�͇���Yf��'uK�Q� �+t�3=F�^Xc�]⎈7O%�@����"�:���P�*�צ�͔��$D[ʒFm�o>��Mc�c�������ͷ��X2���^��C,G:��J;�D��00z�ĕ�4#��%rΥt���D�>�`\���X��EA	y&�D�i���VMݲ˰y��)aF�4{9e:ُL�Cax��2$�ѱ���hxpN'Oikݛ]�&�UR �I�C���m��Y<ŕ��$��h9���]����,G��HӅ��,����m}�}]
��Ls^�7w8���b�����,��w(��yf�;U4ɷ��k9!�kf�r��WI�hس�
�e�)����7�	7N�r���������؇��$����x� ��/.Z
�:�,a�A����]���f��[���_�z�������\w�PbU]b���	�+����"�׉t����!pL2�w����L���n��8G�{�"�Ԯ�H�#�z�%UE6�U�z��7�>�t`@Hy�����d|j��".8BDvk*����F�D��e���q��31So�+Y�w�Pwm�6��9�N�1����'x\�ڝ������
�.�s��.�t���g
�E�b~����{�V���>rn�֙����2H7����,��#�����~��M��*�0�]cv�T�Dju��9&	4��g1�n;�+�
�j�:۾Pj��^P�=n����X7֍t<'��R6�K^@f��G'��S@���g�G7C���-IZ���6U��d�Ϥ�K~������B�ު$��������a7���8]չ2���4��hL3�|;?�B������z(��%�t�z��uK�m�ޕ�����u�&�V��80�� �z_�t�͙�
?lZ�l�N�嚘�-EZ}܁�0��Y&717�uO(K�`�V
CpS���6�J�r�9��e�;��� �����+�*,�m��6U
5�A�I�/,���~>j+�n����T@󐩦���E���=���4b�[ߌ�6>���~l��\����/��OD���h���w7�-FgC(yl.s����9[Ƅ�m�u����!P�L	vB5���?�vY��8�ܖ,h���8Se���
�~��ۓ�t�����pC�������Fĥ�~h_O{�S���Y=���WG�i�!���g̃�Q�T����^D�0��p�3_��UF��vE~�6�? �����\\)Wr��7>���TO�Ou]��Ћ����k����o�A������7+��8 ��p��n��S~�G��7j81��f��8�:�U3���d`�._!x����6�PA�)�'�[��Z�D��C�wQ
��tI���]-d�J-=�T��Qn_�à^AO�<���⩨g��"�Y�XƎ�_�A)�L>+�p4�JvĴ��ԕ�1%͠#�$�� ��յA������>�H3��$׷�b�
q�-�O)"Z���-w���`���'߻��Z�ѥV�ԸtU��$ө*ZK��q6|��qguH'KQ��)�^b���l�Τ���i����r�m,J.�#�9����������$�ϼ�q�Q�g�I��ފ�DL�Wp)�`p�/ 'o9���l�ѠG�Rk�	4g��x�G
d�h�Ŗ17�4~h��f� �W=� �Ä�@�:cF?������4�N䑥�GV�O���
J���e-|�7+�=��D�1}����{QN�/�Ȋ��~�^��4Z�Զ0g�%��'8�0�j�	ĻFl�
D�ӗU�醭=L�� �j���8k������2
��A4��>�am�] �]�|��S��&��)`G��#��U$��	��3�d�Y�N<�����>����|��;��q\"aZW��C����	��a�?KS�%�~����o��.�	��oA=-Qr\M��A�����۫A�ɰ�гQ�:J�'��B�*�e �(���Qvc��@+ۑ�A\ą�p�]d>��/���;9ŀx��)����ms��"4q'_���I��D,]���xn�eC�Ym�?M	?�<uF�%׽�dt2�|����JT՚�H�)���7��Ɛ)��i鴮��ii�'
á/QƭL]^i��|��ά�������',L�s�e�<�����} �pu2�QHXD��T�iAB�m��� �){p�9t,�U����<�\���l㺞F��C�ɝطٻ��W���t��c�(O
ԓ�����.��J�õI�����c�aq{�%5�?p�+��|c�\RoC1����8V�݁��t|��~H��޼ Zn���%L���X�]q�3�4�ɋ���?sNA�� M{�u�=��r��ʷ$�;qG;�g"z����vlʄ�iX�8k4[7��J�<o/�.��޵ ++�sw���e���o� K�/�G�1�A�g�Nv��`&�c��C"���j�t�z�QW1�q����"1�pj�ʄ��i7��litx��v�?�`�|�]�%����X���M��~u:$��d�]yα>���	��b3���F��zx>(��:���H�f��͞/��X>� �l�,"X���H����L��;jKI�s�D�E9�8U�~	��݌'���H���J\@��V{�K�A�b"�1/!�1�e-��MO�Ձ��{��`@�:�-;�P��}���N/�>�H�_�J- ��N�Y��^޸�).����%�-e���8�X��U�[��=\�B!4�!�o��La���0�X�����\ ��;���_�<:wzZ�C`I.���i�V�����*��-I_Ǟ�ˎ� ��<օ��O*5�x���rh^Nk,}��o5�Pz������KL.o�'o3GP��*���Z��z�UV&V"~Z�������CiGsj����.��b~�?��y�.�ե@ق{�ӷ�z���HM~G�����Ƀ�a��K"�;ٿ<<��	���ן�mIFkW�la���S2+�f�]�J�9���3$٤E��;]�|5��o2�n��;��%���IH��g���m?eG��8@�b�q��=�\�=�oE��H���xi�C�<��cf�nS�ڸ&�u����ܱ�O>n����)cUͱT��Ki�2/W�C�#�q�5�e�l%�dK�,���2P6�0���zK�"ʅ�ka�DaVZ��-Mӌ���{[�o9f���a4M/M��$��&� r�C�O�w��������ނx� ���^��`�FE�D6�oVo#}s:b�S�5q�qpCp|!E{���ov��3�ݢ#��o=��D4MA9%�/n�g������?4�!��k�T� 9�������/ͩЎ�	��-XFaJ'��l���������>�ҍ����?��'�*w�b�{~=�l2n#XYi6V#�n�wh~���Ǫ�u?��Dҡ��?��������,%��S�>���~;��VԆ�0M�`p|}e�T���U[`��`ڳ_j�A�zC�� �f|�)J��Xd�.U[�:ʀ(��/}�
�a�߆M�<�x�d1��5K����g����)_N�Pcd��C���q)��/zR��U�z�0h��Y�����߻,�БsX*/B�t�0~^�<�W}�*G�#�?x#�/ݼ:��iE�zi��L�l��;�y��,�!�����yL齙����g.�[�S�c�r�k	�T^U��
�*�<�<=�uL���1�3���iZ�M>a�+ ���A������?��ؑ�n �L�%�w^���F!�%ӽ��k"_��x��z�'�����ķ����2�6ἄX�Q���FB��Q�O���=ڝMn'��K}���cR�Օ�A��H8�%S�'�U���[Dh,�H���D�Bq�1y����'z��<��ME�j��MԿ��Ԩ����D� �B��z�̧������f�S�e�t� ^���{[ob�!�o�"f���	�S�g�Q��l���Hp�f�� u��w�����R�I��=5��d�tR���E��C�ax��	�ZXj��u�9��@��Y�\�W"3)W����{��*ǔ�j�B1���59[��;�j�bˈ��8�x�"�s���Ȼ;VzJ�� y?�M�fq� �&�}���;Z�]�T\|GX��T�Ϛ�|��HN����mg�u�G���_�㱀[:�l��)���juP"ߟA�A�$iƻ�.I�-�0Kx)����s��r�$d4�u.�W~�[�r�L�n��^
�|Nދ��+f57p+����f~aU���a���g{ɻr��9!s�Fh���*%*	f��}�d;��p��O���BxF�Ƕ��!���h�3GDB3ф��nl��d�R{R�v���)<�S�a�Z�����<��F�?<:��+���	R0t�Q'[����	`*ES|i#�ZV&��%�mH��;ۑ۩;�L
k�f���΢L�������[|h�˺���Ȧ�M(z�Nб�k��w4�8(W�MWR�"X����9�.y���*���Yn?���b%�)U�-+#��٧�:I�i`+Ô���{���
U�`Oƺ���<�z\j��P�ڃ-|��g�� �~��,ՀPDB�-�,ʴ�>ՄؓJ��Z�v�{�G+a�I�̤�W2���&Z�Z�jR,n?H��h����Mw�iyB�FT���$�Y`�nZ�l�Jء���n�bb���~�!�b���&y�4�8����{d�Sj���M� ^Fߴ��Ѥ۱�"6R������8��SD��:��W4���~�r�Ncz{��n�J�d��<H����b\	�x̾a��+�~<C�fQ���cѤe��ut���a'ʂ�1s��yy�nA�A?���vX��+B�.�4�b�ZXgM��	�2���ac�M��Q��(ք���~0��.�Le�"��u*$	'rbz�'�ߚ���&_����iv���"$�u������7�V�*���^c@]�|��XÅ2�F҄��]�Qس	4�R�oa�O����c`g;! �U����]�8��T��r��ҳ�k,`�Z�vl�J���dB�?�6k]�C(��v;��";��N( �C�p�G����rLc>Cd�x�oE��U�v��B���\	=+�F/����� y���o���-�.��7�M\�mi�'�L��|�'�k�d�P{N���j�8t�'Sp3E�ݘ�L�rm�A��s��zB1?� ���/�>��9�3H�����\�2-E��1Ⱜo
�Q�W���������e�8߭>�Z��.�^�R�R�Vкj6+$�F�W����2�z>��?��M���Dٱ�ȡ�Y�ڱ~/��ۑ���oT�3 KS<$���ڕ�;�7I�^ �G:�&cU7c������$2�n��ak����:0�;���}��ѵo�C_��"�9�UO7$ �6��>p)ɺPc���1�(��6�l�N�q��L'�K:YI׉/ �G�Ba�����9�۟�2�_V`s��P@L�)��u�\���g�r 1��h����^E�{�h��v/�FÅ�b�����:�Kv�d�*��塚��7�X���J�3���%bG�ϕI�a�>0��ا���Ӟ��d���~m�3S�9���SL�_��G��R3����&.=ݮB�-�=��F�wKQ�t�]� 3���
��B/��M�	�P�ő�#�-�2[���)��x��x����R�hW ��������y�_Q���� ��~	;�e��t�pۄ�v$t��=��R5�m@�s�ôC׽���j��@���qs�9���-U��6"8@Z6U(]0��
˖$� `��z��f�ʳ'�4���,�p�DBxL9�[�t��R�R��Q߀�ZyK�e�骺>9�y
F�:��\�	7Xc�Xba�Q-�4U�������LԆ��_��`pt����5b��=��(k���� ^�Lm(n�p���*�ȡ�u~�L-�5v1���p�n?����w���j��|m��s��@B&v�pߙ$(|w$�i�m
�O�6K�2�q1�Pf�)Zi1P����&���=�cC���E�d���<���D�_��4�
xJ|v��� z��1UQ�n�!	,�����ʂ�TB��Յ�Cܴ̄�\��+PtJG�UR4�� Cvւa�l�9Ҿv|o�5����A*��O��*\����A?f2s[1,y3��^:�����;+�!�,�j�0{�[\ƧC������A���Z�jV��PRJAɟ������.������������r����S���._I��pm�dӏ�2��CyD���p3`���o�$���BkN��[�lf���썜���<@Ϩ�9O8�����Qj��V]�?���#�'��Jz�2Xm([�Hd��.%ɂ,W���K6����A��?6w`^�Cd���X�9�܍�F���|��Jg�>�(�	��LP� %7�kwZ�& �%�nK���C>�蠻�����)5��5��t��oK���uuZ^/�j�_�P�k�̹��3r���\�#�6J~��d�}��6�+�%����2�����,����w��V$����M׎�B���-��NW��tMN����p�l]~�%a�0�7�i�{C/������O�Hܞ.�H'��ޗc��Y�[����#�@2���i�ٗ����X�>:�m1���̍Vˣ��je����XJ���W��}�*Z���0b�尺cn���������7�$o�����D�z��#��z��[�a�FЍ�w��$��>&�:� ;�]�R���?N�/�1E��W>���W�꽪�|�h�H���s�r/��]��@M��t�f���[�.HL���Cƛ��Q������/�[𷹐]�j��^�JFP���KlK��Uuu�U������@�ڑ,��֙��Zt��v��Ru��>&[{��4)C��G�Oo
se������݁�Q� o#�n����ȶ�D0T-Vv���2t���_�T��=��M����y��FV>�J���G3��WM+S�8��>֤�����j?E:5k��m�v$��x����6�[�"@�}�']�g�G�э��� \l�Yho��=�RU�`��t��R���<7�V��?����O�_�s���Z�$:�<�:�R�����+=���2i�%[ �LPd������A�i��r�A�Z��%�_vHT�!�X��`��B�I�̠���vֽ1��AG�k@�9r�&���u�H�k�& �4tBE�l{�C�,��bfW��G��T[,��[�1�h�߬l� �sV�R^n�e[6>��e)��L��%_pU$�j���ÉmN��#XP&�f��"ϩ��ܖ�Z���-m6(�*��YȮoT��l%������D�� m� 4�D�;Հn��,�<v)O'-:��k*K�"�RU�(� س��a�������Ӽ[r��&�'�t��t��\�6}��t�p�}J柑�v�x_������3Cɪ?=l"u{Z�P7�M�=�l��i +-�c�''˭���P��K�q��qM}8����yچ�����&������0���9��WB�:R�c�r����7�漮#hZl�O�gM�w5��T�-�@x���E��ܼ���84$��=)F�����׺Q�t�!�A�]��]Ò�,������S�{?$4�
�K�6 �ӴJ�oc%���ß�����pܣ_M+J�X?���f���|��%��V���B�~�����=�C����ծ|�!�`����sJ�1C0�HYc&�2���3��F��c쎷�X;7����l�~���(�Ϭ������Yc`	:Ե{����[�����#�d~6[ș�I4�h�ݼ���6޷���q����}�s3IeM}�G�Ka֬K�J��������+��S�y �}0s/��5��=:�*Ice��i�ݔ�C�8i�t'*(E�mػN����wρb�I��v��"R��%v;�|�������لA���T�L�u���p1�p��c�W�����e{�0W�X�.�O�u���c��gS�i<Nj�
���<�B?�]9r��m (��Ô�:'�	)�e<��G3A6�L��]Uq�S����Ǩ�u�am��">6��[����t<��� �_M��+%�ƈ�X㋲2#���I�����
��d���{�v�a�*��f�I�y��ٞXd���)/��pyVȐA\�p�I��o��o�1o�B�����2%W����{PR^}1�����ڭ���%�ŕ��dø��o�#p������L�or�HqG~��_ZM�8b9��FRgD��l5@D<�/�-,I�@p�L�v��l�~#X��t�5h�ȹ*�f�߮GW21��wOWoHo�S��v�*G[����X��Ǣ��a����)�G4>]��<È������=Թ�}��l���ڮ^�	丳
YY`Tn���6�N��]�C�E=��j�R�#A8f'hw�-�rLߦ�t�^�SuD��<��v�\�˝�k�f�}�By�F1xv�F�WG�ϕ�k���Hs��Ğ�>�K�)��֊����op�B�ַ������p�ɩ}����ѫ�e�;��ߡ�ʦjx/���p�m܊�H�I���Ed� E)�G�q��� x����AR��q#W��������b�N'��h� 
.����AaFU���u��k�����o����Ijذꊨ��n���b�~F�\Jp4�]x}C0�������֑LO�Q`"儝4T�����J'#Ɏ�S�����K;Ǎ�w�I�]�k���S=���(]*-�cp��b�pH/��}�qd/p��,�9	���P���=t%5���q�0"��:��T�LzQ��
a�4|�}w�(�D?mo�K��+���
>��3��\��sd�vK\���^,�/
��f��A=�y�B�|_�NMp��n�]+�i�S�h�]�."��5tq��X�z�4Gٮ�ܧUb���*���4B��z�։�"����9g�ד��rZ"WT����t�#��{�q�~����VH[�&���y3"���Ȑ,y�>�����2-7,���\+��|�FF�7&� �/v����ձ�YKQ�y�e�*�K��@����궤),d@A���龃r�����4��,۸@m�x�8=ռL�#�dRR��
J9���$D��e�Ι���ca^S�p�8	���G���~�����q�Q!�U������&]�b������ 3�o=)-Xv�f5}��F�N�� E�i˰�׎g2~�D���<�/�4������ޞ��>_.�K��*5�7�?��Z�	���;�c)�+�G{Γ࿜|���xQ6\j"��x�ri{2t��~{7��jh{4K8�ڙ� �� ���X=��P%��F�F�|�S���r�\3�������G�k����U��<fJ�����@����?��M�}%�?,���P��s(�)�JW�>��F~� �o,	CS������8�����<f���qm�Dren��@d+��afnSn �_IK$e��͑��F�7� ��T���T������*����ޕF�7l����t*���*��Y�����<rغS��P�Df<���\!���ȑىX~��nO�ӽ��ɐ�\?�nIV��J�x�ž"x}MO�#=k�vU#z�)�>�t�#��`!������P"�A��q����SM� ��pu�H���?g|u�Orٍ8�n�_�(D�K�6����wP��[ٜu����[�n������ݯ��tѦ�خ]��Wd�l�A�9��bɏ�t��]1�TM܏*�,�-�a�ag�?W���t}
P��jX�0���z�p]�Q�_��,�1@joҏ�V�YQ����̨x����C�+��:��~��6
c��Xt	�hu\�D�0;
鹣�<=�b[r�H���K,njڼ�����nQ�>[����?����͔+m�_��[�!q�ʽ���i
�O�H8�]��~�G%c@�������6����o�Q�����v������\���o�) Y����iC<mm���crƉ�$��Lա*���4߾�6X��O�!�����H,�-�/�P�o5�D���P�iL0cA��t>py~��yL�a�'h�M�b�_�u�'E]���x!V}�*�����*�Oo��U�,��ꟙP9��AK=C_������]5�j�dۆH���#��3*�p��f�9�G1J돰�r��}+�F�����(U��;������ző3�9?2�D��N��ق�~/�������2�3E��,{ãw�Z���`Z.�>|W'LM}5w��nOY��c��懜��#�R}��O/l+�v vI�6�'�#U$Tb�����!]��?XT��!g,@[N�6��!�F��9�h\.�'��k-���i��	s� K��)�t�"ԭ����E���߰'Bx�,N�u�^۔��ܻ�Ns��������{�ئ��!Цb�����%j���F��d�2 OsɴR�p�\�M8j�p�]`�����Myzr���ѧ�����f��y���t�C�AC0��P��%�s2��L���1�8���I�B�U�l܄7�t%�]��^�f�
)Y�EaeQИ�}����	0ގp FGԭfw�ƚ_a�F�C�3���pP�D����Tpf��3�Qb�����)���v��nz���!1��~�=���@�j��qP����T�����b��v�gL�͕��i��� ~^��e�QV��t!��?��O-5�GN�yTF�aW�R`~�R�+l���;�q��l���t�v(����B�v޻1����V|朙����{],M�/#�_K��OB󚧣]�ZR\j��+�6�	n	� ��w�v�����h��xl�o��0ܗ����M�5��o�vRQ��w�9����ӱ��($�1oX48�����l��?B��y�%��z{(��U�c�&�@�f�ƪ#�j��I�=Y4�d���WV4��"���>~��n}cv�lk��V��J�^�����Ҏ12�G�,���}y �::�tڮ~%���<]���C(2�=5�`AE 
ͬ �&0�$E�vg�]R����[����<�F��8�CJ`���E;���vj謎��!LbBߠ˦*���b?s��PP���fS�����g9_B��/�>˯5nx����K|Mg��7�� Ѻ~3���k
�C��������I�������9��l�<���T��� \�rv�<�H�8Jφ ��̈́4���5�q=��*"��Ʊs5���^�YZ��~�6� ��x��ӈ����};�(��y�C�K.�b���vV�3 *7�)VTtۜ���y.ϒ/�y�#oV	g��u��K��}n���P���Xeh��k@����V]�0��$,��5I^���k0~��Iu���;��^^.�c�P͒����!��~LDG�z�7NJ+9�d��pS��*�j�\{y�8]��Յ}�~��d����rnG����Q��Ɏ�r;_)ꜷL�@p�F'"&���SLY��e*�6?��(;0��4����_����{S���z7�cD+V�6?V�7�F?�]F~�^��	'��p_��/8?7Bg7�,b�{���v�F�V1F�����x����Mm������u�$Q���:��������D>���E�}��u��S,�4)N$tiE- ���w�#��D�!a�M���[t��{���-��Z�%��U ȥ���N�}�
�H�7V�Rq.>6Ml?���2�誊a�V\Y��\�YDW�D�`�Ư<>lդ�P�c[�y���3��i��Os��+m@&��}"F9;��χ��9f���cNᚓ�0Ӟ2�y���F���//���l�&g/w���7.h��}���G��UQ> �j������?��ɼ����oωOE�*à7��S��c�&P;�*�����-�.SS_m��ᔄ0��A*�l�ȏ~�����7��h���s�C�qD�¿ݟ%!]]	�e�M>��8����+�F|��b#�����qҊ���mm�w�-�c�����&d�e��b����g}?�X>ce��I���x��rpZ+i��{��G� ���]u��H)�fK�Y2���a�mQ�[u��?��Ԃ�+�J��v�NY�]��hj'���Ø8@`N�M�a г�$�M�7R�J�\��X��P(I��u���zA��GD��"\��sX��a8@�6|g��~������ؓ�~{ܥ� F��$d���|u�D/�8(�qf໦m�q���d�Y�U���,�n�Y�T��!E?�
���`P�����j��5��s�T�m<��ٮ_$�]�1�?J
��o ��R`n��o�[p��e��Mr�3�����H����kۺ�����Q[+�Y���HJ�zޖ2��~�#
0�	�Y��Ӥ�%��Y�J�*.�k�&t�pZ��6ŕ�{�KIH�I�$��+��D�s���[����O"-���%���M�m��[�;��ܼ��VEt����-ņ�Te����Z���ԥ��D��Ğa��E#�:ԩe�����U�	�IЩ�[,v�Y�S����T���E��	w�K)s�r*�i �=QP��tt��%
gU(�|%��Xdv>��V�H��y�&��d������� Z*�P:-b��*��?���%"ځ"��Y?��p�	��9ʥ(l������w�֘%I< ��G��,�ٝ�����$b�c,�r��g��@�#AzlI�{6߯��v���I�3��W@�9�ؙ���� ��*�*���]�\G�zs���0\5k!A9�v������y�"���Z�*1�G���1l���(ڊBN8���w=��t�6���!6�
z��� A<�̈�P�\J���C^嘹�t�=q���bb��a\�尲*��%�Qb�t��- l�$�(e�����⹏�Qі�)}hm�ୖ�@�_UXyDKX:�����{3utc��\�[_Į;'x��vt�� P�-���{d��r�����)�.UÏ����������煇{���t���6W|eZ���t��"Y�놧�=d7�h���*(��[d�}_mD�o"�C�'��!�I2b��,���*	Y�A���)l�R���?�@�� ��b��:]������]R;�w�=�5 �Ź��~׶���VD�)�M=cYB�b0y��D�Z�~.v��v2X������?����ߞ��v����/PrO����2dʲa#,䚟�"_[v��ʴ�1�t�Ҏ�S�DA�EG)l���D��|��}�WS,÷^	c �!-:j�ߏ�&��93 ��F;��w~O���kb�WB3�s`&��{�]�[[�m��(ݏ��[�Q׳aF�ǈ-�fu�>1���mp��L����� �u���.�Y���x�v	�Ј���י�Pq��ƭ���/O����Vtw���-f�b������i��w��D/=�=9+vo�s����e�횏>Q8F:��Q�K�"�`Ri+�8�p ]TB/!:>X�5 w"��`Y=�p�mT}��$��Y�,�p�y�DS�w6U�JO��%�h@�)KLT�BY�J���C�x�����p�C<��a`T>~�Or��ʶ8�^X��՛4Z���O�A������߾n
����Hڬ�U�(���C)����w�s��_�N�i˴���I���%'��]�$�⢯�����w�z1��6���/#B�s�-���6��ܟ������"��#m0�J+)l:B�3'�/��� �XZhW9������b��ΩD����Ԃ���NS�fa!�;�o����ҙ/������V	�g�ݗ�!���}?�CpcWc��m�U������Ew �㰥bI��<at4J3����8�H��Pa%�9���,�0�Hpq<�P��[���.3P0��gf>��I6D��nU��Yd�q/��B��u|N�ᝆ�_Fſhe�5�3#�����
Y�#~I7	(IG�~t��n{jЎ��Y�/�����kų�,�$��ׄ��6�X��ᚮ8z�[���߳�l�#�7[�VM�؞%��,��!�_��wOt�7&;��t�*��˷�r^GS�ve�s��$�UI)b��[+�>��׋��b
a��QB�ؕ�o�^4x��"�(� }C�F}�v<��!%{/ȁf�����YP�"�meΉkqo�����A�q��m3� CƇ�2E�͓��̫�!��[Ό��0Ut�er�]�`��]RA̿��ߊ`g��4Nd.L�͑B���fe��"Z׆s���jV�8𜼨��ԛ�tR�|�{G���!Ame�B��DO���8%�d3�ȯ���Cx���_G�Z��m��QL��:C��IٌjGery&l�m�0��]~�AP/��{W�4�%�@��~k�P�M�ؘx��z>���ʹ��ʀ�|�|�Ž|�_�Y�_'���,U������U���2X�p��q^��2��@�5M�\H�ω�Y%�8SbZ�R��!{�i.���?3�A�=C��p�L�ю�cN~�V�b��.: �?�Q���s7�8Ο�R�Qx�-?ρSq��_W�O(W��D�w׿�����F���~��%�ۃY�u�ʢ�����FԤ�ȕf��R�2��i�z�������T�p�k�b #7�'t��L���/sUC�~�U��#�s�3��;X��gS�g��Dԣ�c�)'��g�\��;B��{�eBJ���-�E�n�X��M4�=e
�œ/$�A�>?�~�{�P�oЬO�Z��!���g-iS	�)m���L!_�HD�Y����[�e�b�N@O;Ԙ�y����?}t;���p*�\�y�.qsw�1@��J��@<hX5�8%���w\9�J������1B��r(~ʈ���};5�H4�`B�0vC��h5�����+u���l��6|;�G=`�6���67�j}9���3Ώ2�g+����H��01?t&݃Ϡ�%q�>��(���j�G�{w�R��ټ
ZF�V�	Sx�yѬ���p3v�����5�K�f��������(lߖN���h'�y��ޅ�TBdE�ո�g�D�h�F��{,%+�\/�ͦ�'7����r|��G/gY�h��^�Ȫ�/�.D�t4���?% ҟ���!��I�AJ^�`���f2,���+�޴�f�9�5_�=HW���r+�z��h�Pa3�w٬r�\$V�gV^jW�_�����s*��j�˓݃*Ӟ�ց�x�
�$v�����:�	�f�E����u�)��h����"%5~��ٳ����6J_b^ o��)V/���ꁧ�/��/��n��H������h~품��Dc�<#��6�{Z���W<Wi����Yi�Wph%q���/0�Ի0C1�"��N��;!�S"b�ⷹ ����`�h-��G��#�K�Z2����|���_��n[�>Z|���if�CO^�
>6��W�ǒI�V\�S�R.��|^�s��`�Ĵa��>���EVV��@./\o��ZI��u��,({��z�g����5�{�f��^���$/��	8�UOn��I�
�*��_0/��4��xyx3�0��C���B�ft����oY~p�T�8�7�a���f�	��F>y�O_�0$����\ae��Mc)q���b�FS�\~�� w'�a�"}�F�,�;קyG"���mF�J��U��5W�ߚʟ�L� [��������\�ha�"6뽅�׼�u�w3=MYzfln���ѹ�+��-�9?&yԪ��N�2F}I����J�*M��o���F�P��_�(�y��%��wnP�f�R�/,kg,���x�B{Əv+���M��X�W�R�х���qU�w��Ga������Y�'�]캓!�hL��g�D!����^�4'�	�V�$���@��̵T�g^��͊��<��n�jo����eD׼���c�W2���f���f[�/`�G�{W�LxWL�u��N���	����t�m�8GF
k����\��Kr�+����}�`��=����[������;&�V�0��Te���Vk8�uMM���ֵEV:��#>K�_�RIy��ج�6�J������y��A�rPD�COHW�[��+(�
O����g	W�����3�A��[������Xts��vҖ����I����B���T!�s�Җ��:-H.�-}�<_/�%�z��(��v�Be��a:uN=@*��n]��
��/P/����}Q�2f4��.w��Y狇���nʰ|8a�	��W'�^�G��G���i��^�\&������c�N&h,L.��&R�
���!�{͚,��{��{vГ�����|�;�B�|rGGj�Bo��<@]���n�����3d`)��z��Tg�5����Z+W��O4jЄ�ut�c�s�qF�a��+�Tb�c��+�4��2\Xq��B4W�U����8��%�^F~ÿ���WY����g�L�J�$õ�����$m��{���A�X�3G~�@Yt�%��q:þ^p��P����N0 Aw�eG�m����wnCK_!�с��r�j�F07����O:����Y-��U��w��C���������j�"Qg*8���"|�IF�_%-��*3�	7x�F4)깈����:��[��?a�������"�=U��E&�X3��W�]��k�^��=�#�L���Ҍ�̥%h	m�F��	�P��(L<A\+V��h�s�����}�z�|�F�%����O>�)�U�Ic���T�z�..�n�e×x@aL_�)"����;�t����706{X��i)�nS[��
�dSi�S*~fM,�d<�5)s���͸[b�H�6Q�:B����'!���2��֒=�*�|�ʁ��޶�\?�)���:}���Vz�C��M`}�l�-���i5�j�.=�"v��	�vv�����\+rt2�u8�>6�u�/��.���ёNӥw���Nr"G��4�TJA�u������0B��9�	ި󁠠8����C�<W�~�q�2����N�D����_��t�5��c�~���,O�3��q3'1&D<)�����h+�݁� � C�4�;�]���;6��e0�`$9lx2&ў��ε򞓂�f��X��� $>��º��V�|s@O;���������${��-]JN^X0��
���+3��$Ob���r"Z+aD�zG�D�#�t�b(aU���Pm�����HHA�G�.>�ap̚	{�1 ����OM� �-^*�i��Vrb���/��~��h�H$e��O�L�G��i�#TjQ��df#�{;��t����"���7\1S�X�%���Jg p5�4��u�E�W ���DN�Cx����zk�hFL�mU�����26�{�ո �u�~k���]{����������ٱ�0.��X\K)�����
T������6\�����o`ʃ�
�{�ߎFm}����t$)��f�i��<��lv�wmE�3k��>�w�ʀ6���ƕ7���@�����b'Rs��GD�x5e��W�l���W��FMK��	���Y�vcOJ��#��:�#m�|y�j"1Kx���e�a���8Ϝ}P�{w�غ��T��2,�"���Z�,-K���@����\
��X\�$*Svi	l��pcA����8��t��BYE������F����	�F�b�a�廓%c�d$��'��=fo-
U�T 1U�vEC�5.n{�p#�9`��$�_����}կ5�|̎"��	t� ���&v�I�[y��cFB�G��h�Gǰ����ZC����]���ݴ#=���\h��G�m�U�X���3|��M���Z�����\Ij��Sؙ0:vo�j�L	r'�N �^�ې0i���=�%�b�*���EkUis8Jl
`�F:]a�h�G'�R��:E2�I�`\�yl*�!�Oߊ�˪�����?��V�v���`%�����z6��&���q��)����t6�C/"��\���+N8� /117��l��(��!ߘ��n06\Ѵ�����Y<�q6��R���� �U��~�k��$�d��@����W,�
����m�/�Ԥ�I��5T���פYu�_��4"���b�ȃD�pړz#�-�&.����B�!Ɗ���*�K%*��%�΂yȥ[�)�,Yڢ9(&��,�:��3o6-�_������=j��E .��bE]GE���V)�gEʕ�G{�lY�e�y���券T������)}��6$z��c:�� ��L��Ʊ*6"���@�Rx.G��R|���`i���Q�u������C�w�T̜O!M�D`;4ٟ�y�fd!�F3�_�ϝ,�q	V��Vn�h�!�ʔK�9 C�Yl����ƒ8ߣ��6���c=�Q�!B�6�I�,	?��'9�C�K&N�"����F?cz�(�=-�m�B�*T|�VشXi����b)��S�T�-�f����������W̫�A��&�5Pڦ̇���J�c�)ӱ	�뢾*G�d�2�f�O�d���[�ÅQP�	(LY�c#NT�g�Y3���D���a���0U?M���f�:�-K�-Ǧ�&�!SD�1�[���1���ӊe��ӷz�ˋ�yNQ��:N����D�ϳ�W�	��t��m���$�ۇ9ɫ�7	sOgT�"�2#$_���e��8���vo���������"��*��@;�2���7P�'�fW��m� Y5�>�s���J_o_a��N� ��j�j�P0g��btr��>���r���W4��&�p��oL�S	�}�cYѳKԛM��>�kMIv�h�6���ԑ�T�mB�WÐ�M{I��Ko]!��'ga��=�Ŷ��ʬ�! ��P)O=��;pc�����mv�O8��=h5N+e2)ϟ�{`"�p ��I����ʈ� ^�j9����HG4il��3�p?(�j3�G5��Z.�Y7�<�����9�v=K��f��n�RKn�{�D��+6��X��#�u�o1m�p�#�Nm�g�8ƻ��d�(�4=�Ӷ��Wo]蠟���ם�{���dP���f./Bg��P�4��NG�[�>,���L�I�i�]ZB�?z��f���u��8q5�������
E9Vk�\��c�\e�	�{�J��b�l#H�a<��z�ߨ�o�CD}Y�MJ�
[1�M|�Jc҃��ϓ*f\̱�解EY�>!��p��#H������$��$��1����1�Q�\�y"rM����+�]D�U2ؿu�k�o͡�r��Lu���[Т&5�3��nʑÈc���d�=
�W!D�ި���d
c�?�&����-�f��(��В5mJ+����Kdx��G\��R���kY'p���	�:����j@j��$wJ:&�����F@�*Tv`�ѳp�Eѩ����8gE��]���^0"������SЌ��=j��!k�=*����yC%!�f��RJ?M�Z1���Svrp��EQP���2@�:�s�1�6q���
��'|�;C�[�TK@����d����"c��Yh�_O"����'2S���`�1�<���rT}c�}��Ai}�Uf�"���/� �T�C�/V0�w{���� �%-Q�9E
Mϰ�j���Ɍ���P�U1��K�qc�y_e���@���x�
���$&H'�񑫁�Uj�d�*׏�yh��2���<JV�#F)	���C}x�广���Ss�D���� ���$������tpɈF��'����|�(��6�Bd�41�s��GcEm��d��P�g�9>�E������Қ���mpv&�M(��Q���iϛ�ş�δ{I����Jd)�7og^�ϟ��,��x��Y�?(�$u���(�����������B�k.E��	р]��м���`���3���!?������|�	��T���� .�ʈ�x�&�+�js\�K�8/�:����Q0?����Z�-oh.��n0#S����ii��1�*-�3���!�kt�t�0WD���&�Cx�Sh��b-�@aP��^��#K�x,�^�+����� ?nJ�H��!���$Is�<tՈ�s��^v9�Ο�θ�dRd����e��/�l�#؋q8@�A�nf0[g�p��Ȇ{�A\�j�bR�#\��U-�Ԭ�����i���bu,���J߬�f<|�'P��$6��G�w��J��^"�双LA�!<��y��>f�=��!	2E�����WiWm��TQ)�-��8�4F�LHX�v�{���5���YJ�H-6��m<N�X�X3�"�[c�'�b�b-oB���j0%W�7Ł�<��ޖ�8N+��<aP���wZ�Ge~r�G1��@�������fˍ��4�]M�
��"�_�.	9�v_�ol2S��lw�C�_d�v�/�S�����r�l؟l`L/��"t�aDm��ヾ}A�z���2#@u��ט_�\�[H���R�_N�K�l_}�=�6�L��Ã#*7�L��w{�h�fd���!d��M��X\��c*�����0צ�X��φ�i���*�3���?@y�kJ�b�T���bgk��7���|Rd�oF�d�?X����8�*8�@�q�8K	�%�)�J�Dk�9$��f��Oc�-�r�\��YQ��7e���#y%O�@�R��(��q�?%�PM�+j�Rv�c����Pzb�c�A���ʦ�W����{��&Xh�;qɮ�Y?3/ ���Ğ���0������Sʯ�_@x���a��2�󧇷^CH�;�[���4O�
��xi�������Fh~����g^0~��� �����e=v��ف�0�6܊�<pUm3�j"�Ss�܃�����/�Y�����У�3�^�����i��?��ue�ل���ȘQ�9�x���Ӄ�1��`(x���L�imŐvP"[�Ӷ�p�ػy�u��$>*+4�H�NZ���@��7~f���!���3�%_�
F)�:���{^��O�L�A,���&�n��0 ��6h���ؙ�Ll�`E
��?x�+I��uU��{����Ȍ�I����]\xX
�,�(�CQ<�ȃ<3�1�����OT���2in7�R�k����":<!mLG>�YV��k�q�ؑ��3� e٪�Z�YT8�YS��1e`���.B[�ŝ�9��FU�ZS��5��L1,�}PW_�ވ��Y�ʳS��&�������[V_��q�D�d]����Z������ݪ�B� ��`���9�I�ae XBm�SE���\_,�����E�0|ӥDS��[�
�����P����(��� Ӭ�_P��O �pW�q��2m����
`f���/�+/Pq�l�oΥ(y*�������	4�b�c��c"��V�//�<�0�|.����'�Ϥ�aV<�m�t�5QD݇suWU.�?�:i��+�IY�Jh+��� |�xO�xR��+A�����@�(�=����"�>��FV�`S��ǳ7�������`Feu�*w�������)&��?M��0�7֛��������Pqmʯ/�}�x]�[�v��PP���m���ybw�7�_M������m �n}+��It�����W홨�������e�?�&:B�P<�e[���� oF�����rM"B�%��>�+e�8�/�o�U������g�.<ez�����U�aKF��.'�	Wf�S���ٱ����������>�M"�VS+�oԵ���4�R�f!���y|��b
*w��{�>��¬��r��Z��=�j���^��0�sYDX���Mq����aq���Fs?9{��bLcp֒��L�7K�iU!�	�~[�*�����.�Y�<��=z�!ZR���;�-��BI���L;l���o����I!�UW̩P1�a^�����W���r*�q��@�Կ�i�o#۽<,��e~&?�}�X`�j2F>� �E���S������dLʫh���zX�����x�P��X*M����W�t)���{~��,`�ā����Ͷ���R��)u�eXj����� �A3�Hk|���w�O&N֛T"�Ȯ 7��W9`l�/!o� ��!�04*���sB�F�Ꚑ�*~�:'5�Yh�$y� �-s�魳6�7u�b�C�P�n����5��Wy�y[h�@�����EOluz7սS}��OYz�뺜_�<��K+��O���@;9d&>���qPu:���Bܣ9�}�w�ɦ�3?�?0?�$��\��o������L����C�r£�u��bf���If5Y�S\����
����x<��3��g,X)f��N���Ƈry�:�0L'�����l��Hn>ۦo��8��pϨ>�(�V��q4~s�4�n�~�E�r@�%�nƦ���0N^!���+�8�����>��������V1��?2�.�����;��;_��щ��񶷝��(kU�% 8a�uyd[�ť*��M|F<���)d*���M�Z���~ׁy�q�jTg)P)��Oޞ?!hx*Y�l��bo�N���@�kw%�O\��տ_��@�הگ@�+���F��O^,��/�7�[R;:�!��P\�Ω�ɕK�P�T�2h`�h}Y2�x1�J612�v*��sh%Z%�F�a�R����!َ��>l䃾�>Ό�5TWl�Ё��po�a=ɹ���	<Er[��yI�r+��\<Z��0��S����$�=�׶)Y����;��1����2&�q�N�����І+J{S��6��$%|�亯��sP f?@�>X�d�.9U՟�����P�x�V��0 �A�; ��ّ����&(����NP�b��&Û/�8c��D�I~�q!(�R���s��lp����E�|�we;�����X���I��T7^�<��.���oʮ8�;�8�{\蓣sΚ�}+$ٺh0�z��{�}sj�2�Ŷ:k�[������O�H�Bso��Mv>�x�L����W_�W�3��z�����
|F�T�U�%�ee���# ������}^�1�B�����VX��g�zy�j@)����_&98רG�oL�,��z6�3[C��n��D���
f��]�p�9FvD���0>L��ၾ��3��@�-L~<�p�j����O�Ur��l�=��z��E�������w ƈ�Z�^!�^���a�EX� |$����;o�#��p��w))������w8|�ؙ`�M�Bٓ�A��Ce��
W��TBW�mW�{�ҿoL��:�3_r뀓g`	�_��5D�����XFs"��i�0�M��Q��(�Չ���Ƴ-&� �M_ϑA�,hv
^��'Uh+W�y�ѿW@p�0�k������+Z^N�!���d��<O�q�3Ц�e5�=A	*��y_)�.�\a�XB�:�dc��B#HU칔�vd�Q�r�*SmUj��5l]�#�HJ���m���x(pQ��4]�?����8(y�vlZ���V�Қc0=�����l�1`-2�
� ��{��%�l�~�����x3�mq��+`ȤV���[x(��y��W���D��
�" C��QzM�Y�~����CL5ɨs����l2t�ԲM������@[�g�]�C��a��o��=�9Mmc_y���ln��M�8�4Ũz��qbP��8a��N� �j��1Jt&I�R�����K쉁��BkJ��3g�-�Ě8�����&���	j���U���a5faRc�A�Q .D���~0�ǭ����񐁹����|-�^l��b�b!����y )�`8V|!y(@��,i��������B
h	J��l~.:���R�l��.��n`gf��&�����K���8���{\c�{�ߒ.o��vY����3�7�]"�v���6�g�+��o���/�����M��&)e.�%Ϲl�~�8�T)�?�*��t�N�+_�4�X�j'���O�g(l]�X���p��$F�YꆄA�2���?E�ZlD6$Ұ�C��'��<�6=f�L.E��	�u5���5c��B���svt����f$�kh�z8��E�|������ċ+���O|�
��D������G�?��2�߻�C�,t��VO�葭T{`Bݛư�k�>�:��v����R5�j�3#���m���a~"�*-d0��At�+��A��{J��������
p����Y�6hx�i� ��&�֍� ���$�^˖��JS�1\� ��+	R�7.����qi��|o���[U��\��E��j<��Wr��l���QZÌVi�8�_�䫆֩RbR|�n��nN�|)5�����Z6T���1������|_��]�6�c-F�K�+l�;gJFY5X��b���^�����&�q����.��`F�	�xd�����y�MU��b�3#���]ے����D�\Y	�FR�����H'	�z�L��V1�~���"X$�!�$\�<ӣH��dD9�i0�5b��[�&_ �J����zs뛱X=�<8L0�B������^;WqD�1A=N�5��X�R'F �����D�0�1�P�;\�㺐��~6���dow��傒e���+�>��[�T���K�/C�q4oH�j�K��qޑ8N	�RPr�6�8M���a��s_�&�.�+����а��M�Aߓ���u/`͛Lf���6zJKS]P`���E�L{��{7�? }5�.�>����&I4�e�Y�r���2�50�]�2����ZV� &������8���t��5V�q�ߣ�*�o�l��s����*1�T��&�(@�zZ	J6s���jc�(%�����]>��:��4� �������~�Rn5���x�4P�!�D.!]Vo(�<���^f~�صۈ�y;M)4��Z�=`��T����>a�}u��H�=3���3j*u�e�mTL������f�"��8�Ϣ�ikU�5I+���L�J���{r8���E{��V���I�I�Sr~e�gf���ƴ>�T�)w�����MtԀ��cgK�p?��nt	���t���	�'�'����'L{�03y�o4E{P����GF��>�c,��6 Ct�_�Hy,������T1mf�V\���W���|�A�$iҿ��Ǝ��2�����;����B�u3▯�M���R�%��*+��ěsn�	c���O�	�a��ywv��q�L��.�@u��1�["�T}���0��*Y�㯛H�5��d|oA�����P�3�Mwi/�����ފ��	U���C�ɈS/��|>K�Frֲ&j��/���^Q�qF�I��w}V����$����U���飛��=f#�_����jPօ(����8=�߀�&�A�Al:7�Ě��;&�Z��VfO��51l}n��ؗ�[���`�y�x�A�^'�����<�����2N�?%��B�����G�6/�4�����s������=v�Cw�ϔ3�I���N�[G�����C��*��R��%�I.H`�\�_[�j�t`W�z�+�awyY�I���&5�(�jl�T�I���jr{[d6���^m���4���37j�A\�'.Տ�#�q�8m+�쵨ޒ�J���ä/��r�ַ�~w&�<���>GB�N��*<�B9��S^����c�Gm�v���НbF!���u����5�O��+��H������q�W�U�d���	'���T�=+E��6�C-d'�V!��S�q�
'F��D�@�vz�	��K� ?���_����oxi����6���ܓI�J�T�X�L��s5��%���d��r�1�Σ2�t����y��h`��j�O��U|Y�7��>�>i�Q��v�-,�J%�Rj��M�B�+ʗ#���Bˑ"�Z~M���	��:Ú�YG�H�Ml�1۠�����6�w��8����M�n�旀+J�K4������i�܁���8KtZ�U�!�kS�e�`�x��	�4ˤ��� ���6�>y{N�J>Z�Z�Xݘ���oᏴ٩�TQ6!ì����0�)ڹ���+�7�|��	iS�ٰ���Rc��FNGU����Gy5��㹝�����I��É����+.�ę�d7�^����q�2�q5]�y��8��Dh��E�C�$b�R�,+TQ3��[$Az[w>��A�x���q��x���>ő��Kjݨ�~w����`�I��'�0�2�G��i¨7�yPa�~Q�&@�<f3�xȽ��YB���"W�6���L��g����X�|I��ə-L��]*{�E-�N�E��'��;��^��7Fԕ�����[�R$�w7�%��2�k4�v�?PЉ�Е#�@��gD{͏=��e���0�3�����<&!.���ڣ�Og0�4��d H܍t2�6���b�9�	���9�9"����zrctM�M�D�(K�z�,��K���,-[a������W��Қ�C,W�����(�@�l�+�<w׵�q�Do�>k�� ��q��=�q$j������X�~ts�џ��������������������
���Y�'k�m'�t?�1����K�hj�*�͏e��!A���(�j�	����
qI�	ݭ�=�v�?�~�{�K>N��/$;Y�mf4s��{��{e�G�a�0��V�sKg%+Y��σ[4p��sc���Wqȣ	CpR�_?]�(���xL��s���d�b���E�r�Y��t.�)y]�FlZ{�;K���<@hg̃/E�+5�ю�噭��m֒����짽�@嫟<S�����3�{�/X#���f�(zI���n���VY�ģ£�`�k�6^�)��d��<Dy�;��Ӳ���[ �Jp�K>yn�*��.��_�6�����*�[�U�b7�VN
���8O�4,��P9��>��ȇ�:a5�"�
����4�v��ϓ�A���U���EG�{F�}u����k���M7��1nB�4�8�*��R�����N��~�ϭ��S�I����<��M@ �1Q��UHtv���4�[��	VE^!��	Q?����0i2�*2�)MK!��f��b��a�V��#���|U����a��O=�X��CD!���i���;U,�&���7S���I���oꑻE)9{�� ^�O���4	�Y���z�K�KmC�=��������nU�dy��Fs���ǋ�4�,� j��6oH�dFk�Zs��G��_w鵅�u����N�a���=��{���[��X3:�H�F���䡔�J0� a�l���-��7z�ex�U_:@}��/،8x箼�ت	]�"e���	<5�\��N��U���:G+��dl���I^�F#�n��q�u&�+�����;-�B�t��Qz�^�ȗ�t�ٛ;�U4Y�x�%�0OU�R.�1U���<2�Ȟv�#x��7'f�B�sz��0K�|3��؂Pk���c6��c	>FuM���O!,�2�p<Z5�v��v�F���K��N��؁A�X��A�2��|�zW_��D�/%Kr�AT�V��U��V�� ����2ãA�������`K�nѥG*�K��Ο�ef��Õe $U���	}6�G�Ƌ���JADb�ta����~4�M*&4��(|ⓣ�;,U�䅡�.��C�KjF���y(�7���������5���=�3�>�Z�%�>r���� �$�ǐzr�
 �-j.�<���/sL�ۥ9NA�knt���k���<) Y�x�HVofR�R�NZ�H�f�0��Ѫ�Q���ª'&��l���Kѕ=�`�8��l��@t�U�1J����x�sP�3-�x��"*x{����.y�`��' 5l� �*Vtg8<
�յW+�q�ٳ�9%�p�;�0����ye�d�C����絏)���!�J��6�	]��k7à�?�!S��ez��%T��XLcJ�H P'�l.@fy�zts��Sk�Ɉ{ez�x^��A}�	����D�v1;���Aw�2��"�O����5��ƍ��4[��A�.���e,��O.��C����'uݒ��%�����޸��|<�BZ�}��_��#��%�� RE��K�Q�����1E�*�Q�a���K�0�o��|��ɽ=�2VҎ��,-(P��t���d�މ�����E~5$���1�ȼ��uL�^�=U��9k@e��1ӂ��eu,mT@t�6�*��G��q���_P��<8[∄-W.+?�����X�A��o=�ۃGe'E������#�n���:��FԹV,*����do���0l?诎�g����w_-�-8�8kB�Rz�.��l��IPk��XHrPl���=��(�-��=�RT��lL� Ip~�S���Oe�X���̻j&D�����Tt���fɌ�E�X��Ҧ�� ?8��iS���_�^��O#Ǖ�_X����(nj>r�V{o3�[�#�Kq)���X}���1Z�E�A�.K����-��BWdl�.�_���'!_�S&���w�qV���9���\�D��᎔$�3m�SB�XB����`3�ドY�z�ma��jw��9�_D�ub'Gu���	�<af�ϳ�b(2�T��]��Ҙ
����e�3�Z�=����:x߲����B��G4t�*HVɂ��6ޢT���Ly%�S���Y���f{M=,@�I�Z�����H"��$�����sx�O"�U:��b�+��d�e&{=Y���#��BC?��?ϧ�-hopb�F
���'ٚPO�0:b�;&I�B�
���q� �n���=&s��>��hބ��Sf������`�W�׬
���2-,E23�>�4�	��9�abARVG֫5�ӭ��kHa9�T���\�V~�w
O�^�c�]8��xm��eS>��M��f��w�bW�l��02j`Y�x�Zu�<���Ҡ��頹[~���O�isc E7�?r9�z���l%�o����y�� ,ݬIѪYޢD`��2�J-Ӷ��g�F���4rE�#�:-�w������[�.�վ�RΨ�#_��2!�[��Ϭj@�R���� ��=4�}(,��K��g܌y�T���@�Q��<��ܤ;v��ۉ����%���1�u���.���'c�8Э�燏3�O��K�[�C�
�����2���vY�|���	z
���� ��:�p��Ԅ�
���Ao���K�̶Ù^l!D�B�0e�Ĭ~���2�'�W��=Q�ݴI� �c�ۃ��o��uI�][�G�Иª�qcO�Dech�m�}Uʒ����$C��=�W�$T'7��ҝk�`Oe���%K�,�fi�Y=�d��������P�Z�p�;c|z��j��kWeoY��fb�&���F��.+�O]H)�`�����8c��ܯ�n��l3�E��o�r�4 ��Ÿ��\�u��\���Z�k؎H'!�=�8�j`��9�:�YP���)[3��
\�ʣθ14s۝F�	��I���G�z!�`���'T�������r���4�x��(G�b���M�(���Gh�Ic�� �,�|���6��朚	��N�g�R2���T�\D	�U��k���� +#Vr�v�DU�[䞧U��x�:G-%�8��S��������*� �oQ�J�F�3��+�1�>��'�Z�H�'EI����v��&���?��$oꌄ�ΐW�u;���
Ifk�-�&�m���U6�"'��`�7b��0�,$�3;�&fPOn�km߁��|�Z*/�����bԸ�y>�!dS�M�@�#̓��x��4V��䑲n��k2y�fw�`no^�8��;آ��-����\%����&EA>�� Ǎ/�D=���9�"{��W���sUU� �<�S�_�4!��N����0\`���o*��׈.̓��C��$��BϦ���H:�ڎļy}�¯�Iܿ�ʃ��z"�7Ǥ����lA�?�o�{@�sb��
�%�+e�]�, cbÈ� kT.>;[����OsX���c8>>��R,��7 u�q�O	v��m�=G� �&�#�&���ȸ�ˢ���GǾ{��-���iq�J���hQB�c�T�d��E�����
\vE�G:7�d���i���4���{�tP~ke�̞�_[B���KATZ��L�;�ڛ�QJ�K�w�X��h�/�׊�(�۪%^Ů�o�����%���K|ZgU�����!���e�Y��4���
���/���V���M�"�8�W�~t�ϔ9�~��˖�L���
�w>��xkB��:�}�l 	�t����qGjv���#��o)-�O���p(�3�+)�w�|��a�w�q�����-x���Mw��'t�$
��r!g��GF�X̏D�Y��Z�ڛ��<�x��g)e{����R��ݑ	ei7S��gE�S=J��b��*��G�֨���E4���v	�C�!���k� ��3ɩ�����e�Y�E�&�0[t��#�%.x��w�;�NPd$�<�vt3�5N��-T�����ñ,��Gy��h�ݭ��˵I�K�������H>���
�q鷾z'G�)i�`�V�h\i��B�5��H�C��p?��u]�b��^��.�����c$eE��7nl����Vb�u���6Tϒ�G��pXΝ%�Vl��x�������Iɷ����� J�K�"p܁WB������ sC����2��  �S��#d�2~��"� �e��;�Hv�Z�i���7P=���oI:
�:!����a[*IBr1A�8��j��i׀�"K�5��!q�.�Ʉ���l�����<pJ'f�^����>% ��v�h��<G��(��11Z���p[�R� ֤�~}t/�5�����@F?>�N��p��\�Ĳ�Gc��D��0}V���Ml�ګ%���&���B�����������h�X�������y�x{X�ϼq�s����n[�Oa�fa%@�g�KI,�ލMl:�:�j2Ք�+=�)� L��}���$ם� ��Æ����W�\����*�qaiqw�)(���bTRj��uPTTq�f�f{��V��Y�10i��p!1��oY����E��>)�.�&o����l��I;M�b*�E��hD�{/[k�����%����]Xw*���eI�P���=�^Bd�r�8���̛,�=���O�[�k��j��Y��v$��� �sM<z$CaQ�.�1�9�_����CPJj�6ff��-v2�)	��)�D%�Ck?��� ɐ�� ���v
pЪ�MEP�g�Sq�sF;%�ޗ7��`��8~��p��B��lo��]����o��������k��+D����c��|��Iޔ�[+��0ƼA-/x\�6m 1���*#��E�w���ܰ:�}��-���V�ue��r�I�a�ݝf}�����mu��ꍶt���ن�
�?dM�������i�´�AB�6�[P�]%�^%V�cu��h�
�9�ɻ�%"�0W�
��Q�;/������i#��g�����dUH|��q���;��j{E�Ƥ��;�<C�N�R �8�s	ߠ�D6�ȉr��o�d�D;e�q\1�Z3���דGPPx�ŝ}��o#`dx���o���I�G��(��1���[���3l�!��.Wr7cFo|21|M�������̓�`h��yU�l���&-ުϨ�0���v�Λ���\�lt8iF����p��
Z�������?���:*"�Ol,l�%Wi����Ն0�I3cEX���Q�D�A1�<M���.����c8!�}�P�A:�w��_�Tj���蹘 ����L��P�p��n9�6�����A�6^v9ӗy���ע������~u�}�Pū���N�/�jg&[�s���:
&�Ӎ���?���3Fe6��v	ͧ}ʯ�jN#�Q�Y��'N�<�'	cڠ����-�H-��@��y�/�ٕB]y6�^A�l�y �~鈃ng��RB*9!ꢇA���x���}�f�ĉ�Z8���+�AJD����v�*�{���	�Y��i��T( /a�Z�#��<�T1�K68T��R��t��L��Ȳ�D�
��CQ��7���J��]�rjKRݕ?�^E��.�R�����<��j�����6��*��R`Kw��iS\y�h�S9���*�os����w��E[�˾P�	�'I�R��yge4�e��e�����o����4V!�)�k
)�����X�2ȴ\�@5u�� IF �?vyi$}��i�B ��z��
�=Vf8��7a��p=0���_u�� \����:a�-vڒzZ8?��]�AUF��v%�އ��9A�o>Fuڱw�!j���ȣ3�'����r�1�7������u� ���=b�����g�0�P�1L�g��,�n��X����t[�!GUY_�E5�ߢP�/�����GYH�W�ʡ�?T;"Ι.�6��cn7�.�w�ַ*����f�|!T-� �L�4e4��.��ǩ�> *�M="!�a�hD�5�k�[n"�Kn���k�FD�hY� ?;e��ds)�d��Oa�7���*��>@0NN5lʬU�E�0B��T=Gݕ��w5��Z���H���7X��t�Ķ��ڥ�r	2h��w���,���vo���<��G��4اv�ƗG���%8y��lQ��8�I�+�3�N�כYX$�7e�av�����$�}�0 �í7R[t�@S�ՄsS�f���P�ep�� M,�.'��5 ��q�1)�[Yǉ�����q2���$�E	<i��tEc<l��JN��)L$���O_�ȟ�菱�Ѐ5�F����1�}/E��뵎��Nz�D>�Պ1�&ć�F5}Y���,����%8� %�
�+tPe�x.߮���(A�+��hGn�J%�=�S��[�A��>=�"���&G�&�ǘ��9�f�w�(I����9��'�}<>Iԡ5���XY�_ڲ(6#:Lsߤ���L���	���0����0�*/�sy�@�]?�e���<�P[m�b��ħ"`���_��I9����z1C>p澉H7���Y�ҟL���,��q���Rb�r�_�Ƕ/\q�J�2L"�g�uo���n�F!sk�M��g�Eۤk<�� � ��� ��x��~eth�VV�A��<*h��s��-�@�$����k����
�-Q����	�{��Lz��3��d+�t7�Q��;Ī:�~�������(�ʚ4�h�J�z�D\��N�9w�`v8��:��4���~�K%�pn8`�z1fB��BY����x�X�ɝ[Š��?�����L��$�Ь��id �$N8�憿iu|�V�e̍;�jA�ʛ�s���ΡU� /������g�s���Ĭ`Uʵ>���	��8I��]9d��gp��ahn�r�]A5vS����m�ޟSź0��k�8�k�ȗ�&Q}�aN�:r�HYݧe� E#�,z��J���*����Yc��˸�e[#�ω��Ə�۞@�V`56@�a��R>����-ʸ/�������8�@��z���d�=ӝ�nb�*,w���8����fOrMr�of��}�S��;�8�=���%O����A`��䷂�"�M�G�9�8�	5Kv����c�o�'9�����@P:���͋��~NW-�e�%��ַ���@���z �E��ﰛ�%�{K�m�G�,��5�Bh����>�#݇��w	"�G�7�w�%퍎� ���6�F{�_�P2R��.F���o��=��(��2�{��I�y)o8���!^����9f���x.�DKZ��ܩ	�*�Z�o�=���v����u=���Y2�Չ`�EA �CB3|o���X㹌p�]1���8�	���%�#�]��`�`��o�l�*�`DAu��B[I,���N(��i������j� �}	���"�,cu��_rQn<Zȵ�/!xIAc�p���t7�i<�h`1�5����0R���;j�L���M0
I��O<`#T3�ý���m]Ɖ�������1�-���!�o��e�y�3V���������H�S�Vى,M�n��7 �7-S������ތ< $�c�y@�ؑ5��[����L��y!�)��25�^�
 �[֝1����x�E?�ֲZ���^h�fx����@Jb�����ͩ�/�;B����֩qs��E���b�Ȏ�S��TH��&���;�����ô�b4�q��b�H+L�%��g�oёn�����T��=�>�K*���c��������D: ���m��-6[l�����E{�'^�<" �>�|6K:��̎�Ņ�UxV3=#A��������8�HuPZ�wgYݟ���#:�)��Xt�/�.���r��]U��nE(���)�+�����%!Vt{����Y��D���P����0�y������^���Ko4�/]�/�n)KN�\qǰ�	F#�	K�-d��-��L2���'l���'C�꙰�[S��@O�:r@T�ɨ
cv�D`�E���|���'gk�[:7�Ot�B�>�絖�tG6\zWkL���YT�;�;�V[��3�Y�c�864�m���t�C���܆pV���m�WۓX�K���������
f�����
�GںC��=�C�*gD�%Kárƥ����݃u�Gv��7��v9���7v�ǡބ+�� ������p��-D+�r�~�!�8�������@��QZ� �+�u:$����T`:� ��;�/�d&���Z��Cc�ݣya���k�/����*�4b�y�o����Х�(��n�� 3���'�j7�"{`X1`~��M~����KA,�N
�� �6��	�$����s���JB���ph���5S
��<��Wqj2DT͵����O��o02�=��(��_;;�Ժ��n�����|�U�
IQ�	5��(�Ι#��ԩ�};6:_"VҨ3|�����}ٲ<�{�X��&N�Q�G��P�ό�˽��h�N[i������i���Ba�����eO���2C�_t����@`�(d���tM�Ȭ���#�Q��'r}�F��h����Iw�4̚ԯ�ʩ\������Բgk�.맾�;'�a]%џ;�E���������JԶa��0�c&.�:�����@�4�pJ�̅���F���x~��q�vɉ���M���2� ���G�-t���^�8���^5mrӶ��Yp�l��� _Ԕjl����^���W����5�{n�)T¬�<�[AM��mb5�D�3��^�*�^�W�<��u�/(��8�8���e^�:An�TA�RU�uY�^T��C��awj�+{�0��|�qs�9��ub
��`����D�E�u�X�F#���Dۺ�I�b.ס�6�@��e%A�ӌ8���|���)o��`l�c����n����񧄒�|a�4�5հ!(���]�PY���6�o�D���q�䚴 *�c��:��ӈ�R����cZԺI�{JJ��#޹6�Fp��Q�9Ԕ!_�t��*�<�}詗�UOXMѯ4��1Z��k�?�D$ܗ����(�q]6�Q��c�#��%��V��7Z�(�}&��&Њ��!�����&<�{���־�<Z=��a,�r���jO�c����p�QP?z�����b'ޙy,r%�Xq�,�/��P�!Y2HȚ��=��۳����#���7W�}�ڿ�I-�Q�Չ�708�
&:��p�Hm�t濅��?Tq;�f{3q+'��[���ۺi�W͈��j�e�/ ��Ȕ��gҢ�(Q��5�ݷ<1��0Ue�x�F�^�s��e�/Q��]�i�j���e��Y��Rc��$�1��� %Vl�y������ӱ�T��ѥh��"�Q����It���)Qش��[y1�IQB��#Zl�[��ZE�{ �u��K\g����ϟ�[2���Q�@�%j��N�ʣ-\�B��~�,�3���a{�K�@;j>fG��&W��A��9�&
I�Y1�������5��|��郂%#��V�K�����C#K�+p����:�z��	�W_O�6�H&C� �x���<����@O+ �$� |�QYX,�t��Bk����e=� 9xF7J�����S2
'�N!���N�L�ֆ����0�)c��	֟�4�$�A�'�I��-=�/*�D9M.��X0���#��֦0�I*M�"x���T�P�y�ާ|,ϋ:��>��Tp��0=+WqٻN�S�7>*3��<�H�!�N#Ym�BTLL	^b����_�����j47��{��W�i��[0�ry>� ���1���Ŭ���@y���#�>o��W0�Sɵ�m8]���Bb�&��Z�q�\�`H}L�%��b��*�͢�0���p�&�Hm5SJ�f4ڞ���MR�]s,�qpk���Z�b�H0������w�P�t3�'��l@_�1��fA)��H94�H�%ޫ�2fP�����,k9�@�y%�ܭm~k�f��c1�ٙ5�/����~|lwR`O �ӊ��!?&�'.LSތ��]�=����yPL��{���d')%A�*5��ޔRCΧ�T\۴f�o+���&���uuF~�Y��B��F8�vPAF��(�c�>��_�!<)��^�t &׻ǩY��U^���b�ü�����J"*���������5���C����wRO�	��w�#
����UT!*���1���5�-��<h�,��NB��K��b\�������(D��;dg������q�I �c��i+H��ud��w��*����J��Ƨf�d�P1�q"^�]�>D�.�|���#?��`�h��/���@�l#Cz����F�ĐR/D~{`���@�qF��}N!
.b���&.��(�
�+��L\F�����S�J1�ɧ~�tYi?�U#V=��۔�s)�MB��S�q�R&9�e��FO ǬZ�9�s�3�Q$P��R�$�:��t.��!s���Y�����,|�s�_O�Y�JQ8sq��n��Z�A����R���CN��B��`ݐ��2#E�7�BD�tJ��ʡU{����t���қ۴(��3��q	2W�%l1s�Y&���<yXM���&{4�,1�bӀH�m��D�~��W�I��'�S%A��QZ�狌�r�u�['�oX�hɇ����#�x}����W���g�Z罦-,�C�j��e��~����f��M����p��P
op\3��=�)G? j��7�f�Ԗ5n��
qUl���kW��>Y�=���;�����Њ�o��v�a�[�T>CIw�;�h�e������6�L���4Z���+����ֲ�C�
��y�ţMr\k �s�4	f��#������v�g��ŀ3�P�|��GϏ0l=u��ozչ׸z�m�T|�E�����g)4�$b�U�%8�R>߹�bӸ���p��V�r?��N� B�l��l�7�0U��'���k'���'��w{x�_D�����Y�߀�[�KA�#k�sW��r�x��!S[�[��`ڀ�g�-a����Avv�XW���W4�f `1i���U�~�pA3_����T��0ES�8G�+PZ��t�y�|L��H�!8^�j3�ڦ��"�1UN�j���SY����tD��c��G"RE1iD�����n ���_K���C�B�7/CI_�fUE}+E�f��ws�s�l{��� �H�1��yi��D�Kd����Bn�șp�����f u%��*��@+g�ϊ'�M?�i�"GBb9�/�PKԮ��XTʲq)�Ò�Ô���GO��Yw�t76�`Z^͏����4P"mPqT�b'����b����+��ɄB{^ss\��V�M����#�a�Ir�*v̳�-g��r?dY�XT�^�*�Hf��W%�I�2o��j6�b��OwcB+'���;�^/�S�3S������z������bN�&(�r{�p�V�� ����H:�K{0�j�{�����A0�B7?�q'I��T�J.�yچ���@����7�c���X:u-E�wI�_`Y5��o��L�,���[k�7j���gKܱ����������9��^�Uc���4��	ʹB��/@q֑R��Ijm��25�#��o����æ1ej}�|�����-Ask�Ƅ��y���vy��x����s��ʍϞ��u+<��6R�F<ڍ�	4�JK�+���%�o"�-zVa�uh�W��{���zSϓ�_!��t��ĳ0u ����KgO5_����	���5��QM�_oއ��~7�E+h�D!���O[F�H�~����a�K�!n8z,ۛ�`c�#���a�(E$��])qq��CX��\�M�g�Y6����:�Y�h*�`C��Flrgݗ^L��صN����A\�1O�f;N?$�7]H�pb4�9�``GR��� ��k�t���ƿ�}�O���C�9��ݥQO�şV������9DW)�y��ܳI� C$��+��ic����$U���?�Xu���<��43�,2ӣ�!j>����Ȋ� ?8Ůo�=5�}4hdKPv�^���{\I܏�� ���_=��mR%%Q5fW�=ԫ$3�+n������S���9���'��É�1G�6�Wɴ�pi<u��:���mQ�?���$�{�Z�ad��:�FG��6���r���x��L��F��(s����,�����r噡%�iQ&zs ���c����ID���������r50B�Љ)����#�dm�4`�����
��u/H�p��C��S�(��\�����ؒ����U叴�~f9�\��q�N�����[�Ԧ�K�S����b��w)�āŦ�~�R���H�2�Pz�K)n�li��);��� WY/[���h�e>���3T��9{�L�vĽ��V�� ��Z��ɣ�x��lւ	9�r H@��������~$)�"r�ԧ��5"2��D��/�hmf�ܪ�bt\��B0�,�ݟ1����=�������_��ȫ�`𨔤�7����V�fD��b��|R���$�O��f��ѻ��_`�"2Ϟc؀����\�j؏%�b��>������`x�K����J�6v��/MK������AG�$�z��q�9A��ӵ�G����N��LaI���vY�LpK[��} _f+}��+rv�ċn�L�d�����çQ�c>o7#�zb��c\�8�vW�"pId��e���o���\�� �Y�����?�����:lC�O3;I�pA�$�����%���ק�Z�Ic��o�� ���i��Y�];_J^��+�ߪH���G��R����ɔ'�f�c9-Aw��`�4����!�TDh6�������^��B&���CGk��N?'������-��m4�*�ͬaN@��F�#x�r*�=l���-�h�O{j�F&5�������q��F$8�z{^=x��$�e �챍#]X�a��8����~�����3�84)`yj�D��om�3>�b/�wV�%Fݯb�����%��G?\Ks�fchG�I`U����]u�(1�"��}!U�g|�����c�a�A3<�h;4���sS��)���Z;ڏ"h��&4m|@�"
tuLn�Ҝ�bϗ�I��)�����O�r�_��,�_�xm�&^�����Ov���)�S@�^�u@�N���N=�'�V,��q�>Q'����T���F��0Y&l7s�GF���3[��שA7��4[�vf�Iw�4�A�m��0nx[�X�L>������ʷ�23��*`]v],߶�ք���K�v��.w�my����&#��0�8=Q�+PQ��P��<�B`]0]�=%4��I���,������G#�+���p'�|�o�����
���׬O.�s�&=(B�4�8�Lي}砺�r��D���O�:H����P�l
Y��7��۸��˹�X�� �N��X�͸`j�w���ϖ�?u�r@�!�	RYQ*�~0j9�|����I��Ry(�j�����\����0}]m�IZ�WL�Ys�ڎ�&�z�H��&nB?A�^��UR,Iq�M��.zIy ��뺙��,zD�K���T�?>rE�� �d��z룥V��1QG��Ĥ'{(�B\4)$�9S���^�r�:gc�������l#?�2�'�KU��_%M�jF0��Sn ��	[Vpy��B�b��U)-�L�"m<M��*ȭ���?�e��U�G���5�����/�9W==�I_ԨG�k���i��v�T�[��yw:�Ǭ���ģC�.��A(8����!��wi�{�?~�"	����{�
,��_�����l~�YT�p�<3��!��n�o
B��|׎����/;��l����x4�%�l_;��+�����&dy���q�I��&�����Zw= ��Fj�ܞ�>����mjs@*�<�5L���.��"&T6u;�����D��Y"�"4bG�˨�"�xT`���!$��o��0Dg=��f�yP�$z�[�����\e?�O}e�KK�a:;;��{%t��z���Z�I�[l�����p���͚�0�ֱk��1�����l0	ԁ;4g���� ��S`���� !��&�H0�׈~j����~aT�y7|h�^�3j`���������VH�OIyr )C1�9�I�ǻ듯���R�Rxq,��3]7VT���E*>�x��:��2q2��#�L�0$tH�݈�w����{���ź����W�h������c�+x·�7FݣY�y2�J�oF>���E����5��d��Q�@V+�,�_N�¶���,��8%o�,ó1'q��B
r�!��Gޛ<J4��|����p`����>��j8-3�s�c@Ω���Uw�Ϋ\��\&"[��C��*�k�΅���@3ap	����-F�ԃ�;g�<�܁��9�1�&p���x�+�o�d�ā�F�=u��=_�$�P6A��A(�I�5�J�ҽÕ���;����Ko(�x�Hw:q��6Zqk���o���?fР���U-�-��a������bo{�����w2�;��z������o���)|��Kl"4ɵ!��[�l����d�N���~��򲯣ED�����f,=�k��u�V��5=y��)����9�'X�q���ͻ���]��H�,?�ƶG�h������RN�K�{���������Ln�B[�0e4�){t�S��e7}4��	�QJ%����PW�r�U�q�bw�ˢX�#�V���U�rd�9�a��x)�mc���8��۹�m�����Pfɛu��Iond�����=A��J�Xa;<"�
��a"��3�G�$��LU�������X4�й!]g����p�G��	��8&hsbDW�� >��?+��S�REӨ�F{1GT��Oܲ��Z��G81(�%��Bx����b���1���9�ݮhֹ���1E����%�#u�F��rV�\����dc.ژ�a|�(�Tg��t�a9�ӎh�oc8�1 �m�cj��+��H,�S¦�)��{�M&��u���J���)��ABS'�-L�m`Q�ϪH�(�鰀Z�_Vz7V�2���` �[;��+�O<�!�U<r���5�&Y��e|�-R��;���6#1�l��������1%�:<wG�ѕ5��6�������N�̱Yr��@�?�Ί|�ta �\=�`������0�e|��nAx����0���O�l������v�u�'�ؖ�Z�|�C��Z}�cI{��X\/E��}���5�X�69=!rI����˞�:J{.����8��&��&@�o�s�u�mx
Hґ�蒡��a["�'��V�,P)�
�gv���i����5�Ӹ�L S�j����]n͛Q
,p�FD�v.�$9cK|�Ui��D>�0�0�Fg`�b����b��ߢ���J�ٱ� +\j�Ʊ��Y_�DA�\a|D�Z�L����gY2� L��s��N 6r� ����R8{�D\�^`��F7���֋�Ȃ�6�.����,���e	�_T����`�=�x�3�\���Θ�?A=���He�'�Jw݇1>�WwJ�*0�����W*�&��
R���h���#�
�j�\T��F���y��<4Y�K5�� !3� t��^���
QF��ݷ��G���j��`d���	�+��w�\[�*�GB�~ār��O��KJ�&���u���HB��@����d�#�8�A0�Ӹ�ѧ�� ﮎzX91Xf��8)�?���:P���9f6��Ƈgn���n�;�JJU�ؗ����&m,�!�3T����E�/a�.Q;#�?�E=�_�Eu`7F���wj��ʑ���;^�����e�1z/�X����޹����YG
��h�oFV��K�N�>�����ÃF�/�C��C�b(w���C����C�+�4$ �s7����+�t�,�]�hN�b�s�㓥l�3E�k]+ۆ}�)<ؼ�G�\���Q����Kv7�뉌�E+n*��w�y����՞�*"�X��aI�H��8�ڸ��ՖE�L�<�'$���9�w�� �ޢ����ae�2�"�=&jq��ot�#���k�r	�W�$H�<|����/��<A��"���X����$���?m�8)6��"��6����*��S���)e$@Z�B��b���:W���r&\u
>,��D�`Nk��t�|9��/b�g@8�բ(��)�G�G��T�� ���wA�����J�R\qG��i�z�x�������u��ܫF�a<�N�ϪK���K�h����y�ו�Pk��p&��?�v'h���\��-�0�M,����(`X�I�
9����cf0�t�TY��^�*�n3w(j����.�Y�(�'�@�K(mU������ �2K�%'�T��٩q$)���?Ţ����=87K Y�^�ǲz����pX���ْ�N���"�������7�W�6�[�W��ߌ� y"��s�X 	��OD���ˌ��5k.j��\��x>�D�;V5BA��X�$��3{c��,��Q��N���#�H��Z��E�_l�@LX�ʅ,�z��wT$�\�2��U��l茄1�<)oda�0����z)� _�����\6@��78k9j����_�U]4R��'�ܛ��9l��p�쯗���!�A2�цZt���J@�%`'��i�)���^9M\	��Ŷ{%>��M������^���Ԫ��'G�c�t�)�>�f�8��!�7i��Q`$+�<�it�_�m�gB;�!�j�>bd����7C�XL�M`�i�N� ��P�<�����e�ËS��%2b9�;!>G�t�Ǡ�m�+qx��R��7�^\|J,��U�p+�z��5c��EN��'���G�=�g�H)E����W�8xIY��k��e7�b����;�>K�Z�i:e\�X��<eu�;Z�_NGV��K���k�x1oȟbq�X���?�y�}�`2�Y��E��X�l�ic��f��$��?���G<V�'k���@"`}��u��M�t�����J3O���Ƅa�1��;�Q魧��T ���R���w)��Z8�I.3c�Z�:��jf��h�6뤠��Eg]�JT"��IO�rIp���!KU�O�rP���v��[��U��e��ITT�.2"uo�ï�$�;�R�����+�nץ{"�9�DͱO�C#!X`�;���A�a�k�N�l�н��V@2٫w�\�MН�C3��&��8A��7\F��9s��:��w����1/l���̐��!��w�y�G�^�(Vϋ��fN6l�={F[Q���?7�a�e��������O�.�6@e���;�{J�n�,��O��<��������iq.�
��4<�+#�N���S� �X��g|��� ~�!`viD๏�t�ғ��DL��&$�B�@$��2�Yz�*��|��*����$�0 ��P!P���L�`���Z��R���E5�@�{N���$�{L��_|�M������3�䅮v��� h���y������rl;��U]a��H�W��)m6c��C]6��0+F3{2rgVs��,q��x���U�Ο@k��z�P�%�3C�>��1��E�o X��d�<M=T�����T���lGM����)�ҳ7^1#�CBZ���Ă�T]�:���Z�F��~����F�wcA1�8<���"��tK/�	Iؿk2�@<Y�,�0�J^����	�x4l�V�q)�=���P!?�G�
�Ȱ�c�tv���
�>zss4��I>�`��,5�%#�*���e��%�%9��u�
߮%���Y+�L`�Ud�z B�m�=�%����O �k|�c,q�N�8�#�tZ��l��P��W���105��%�7�]n(M��=��$�sљN�%a�ӳ�����a���О���3E	\��crx���U��U�-�~Yc}0ࣺd3oJ�^������e��tX��7òc�>)v�I��1����b+_'�0���B�xA�����0�u<��q�?����~�ثg� �����B~���|&����]'Z��1���'��lLV� p�5l.��p�
K6P��7���� �/�*�JkI�P�)E�}5��Ch��V[�~�����OʦJ� �ɝ����3����e�ЌPk���3�h�'8u4_�����A����kF�"�]�X	�@f���x�RV�zMO>H꬗�̊����.U+��|k`��J����Y�%�y�]F��۬5y��3�M�ը���졙��9���gؠ�O�;�ǣ�����N%Q�>%�>;�h�O�!�R�5��^�5�_	r��k�wnB+�E�P2��y13����nP:���S�,;�Y;v�f��$��̹���Dr���P0���ҏ�h��'?$R�i�Ǝ���� ���.*�!��X&��!K��2�Q=YS>0����QJ��q	��Ŭdpi�u� ��:�#���|z�lb�ZO�f���k�Ƞ�w����W��fe퇪�^32��c�4"���Ӿ&+c��N!d_bw"��C Bz���s7i�{H���t����ʳ��L�u�y�ј��r�ђ%Y,���r��ؙMwVZ�N��ݩ=rr�=k�7�fN�	X�&}7I�68�{.�c�W�ο:���X_%���.3��!c��wH�M73S��:����$Сg�۬��ᡴ�R��X��NL�Q�D��P�Bu>&"E��~G�:��~ʣc� �Nv�v�+� @�m$�.@c6/I�ґ;�C���([��G�yl�}�9�A�U�+�@!T��AQ����>|Y����&����2z�N.�S��Mmn��?zC=2�b�V��BY�8��	���T�[熏��^�]Y��w���N�O��-hU�P5;;4�!��4|.���%h�/UX�\uΦ�Ȃ����K��ᖁ���0�4<�8����2�W�,��}�������&�%c�´�oȝ�O#5�C�|
XO¶��7j�uthA�[�^Ӥ 1M�ӝjx�ڍ��-)҉�����:����8�k��B/%�ɌxϔMt�|q�u����#2z�g�����-x�7��n��ۆ��V���\�ɓL�u��؏��޺a�<5oX˭Ͽ��yc>W��6��f����m���I�4τl�P�Br^zk	M��Y�vo�n-IpŔJLv�=^���4O�=z���%s����N�Fzj���w����G�@l���BK��l���``�d�#�},oл���\߫��n/�b�D�G��j�n*r�t����l?�ʳ�c�m퇴4�f�&w�y�d}x�^gBh"�,p2��P�	�o�<�ڧ�r�Peˍ�]#��J��Z'}��P�M��U�F��(R�$ orQN�5D�<(;hN?ZDm��gO
ώ��DX�,%1mG���d��DyF�m[Ҋ*���U��`�������:i����>�� ��n�0V	���eX��D�1l���EՁRu�q�l1	C�9�ռ�l���;Qp�R?�3�P`y!/0T�8�j�Q
U��j�â`�p0�����j�ƪ@s�OT����l��;G���H���B]hP35����PR�\e���a�b�3��������/��20hs)8�ps�;�u_�^-���9��e�؀!�F�^�-�k�����8g_��G{7o�'���*3�Si�КpB�u��|KvQȇxJ:yΑ8���&��Ue�h��v�X-����V{8����75kn݀琷O$�{����>����`�]A�����W��+�8��M1]�<o)7��$���aª�C[���|��x������)c�U�_Dj�!
��P�������0َg�ɵ����lM[�����(��&� 9,�a���-��j�TY� ב@�kh���^z���`Q��
I���'h/�	��Y �����Y#z�?��n��y�Z�O2$���lB�.w-���3��8�A`��9���mDh�d�_q{���U{-��KՈ.Ֆ�����U����皁4�7=#�pteWp��O�}�*+x�� Gz�*D	�f@�������앇��~�������n`����d��k����e�T�TX� ̡�h�ձ�[tH�g1Jfx��/Չ3V��y�`bGa�cX�m��fo��j؈	3��$����,�$�=J��+��&��� � ��f��1޴����R���B��9���8�c�R����+�@֥Z����+ji7f7-�u�ɶ�Ρ��(%�(��i�P�AF_�W^��&i`Y���܌@@G���ּW) ���$zT��L�sz
���!$��e��{+d�iJ��A���=z�4������sQ\� �aB	���/	k$��V��h�8��Sc�f�(���,���c)��q�U5��NR�/�:��zM��6(�H�h'5��>����U��!<�pΨ�2~՜F!kT��TQLJ����T��:H��Ig[��q�D����|*4!M'�>xz�H�a���#ب+?�����?}�[Ť�6����*7�}P�\���kc;	r �����$�פ����E��k;��2?u�a����a홍2�Qw��s�Kf�H����^S�a�,?͓n])�;�Y#�
K]�� n�(R�����!�(�Z�G�I�v{�Z���>Φ)2E�A2ʊ~�5�
*ʆ�{e�����.-������ձo��z�]A�?�d�>�̙�gՎ�[��y=cXC&o�w��uEo�moԛ�߿-����΀�M��`����
2��&��mDPvr�'#���S�{��V+�Y�$>hf����A��u����E��βXQ�r�\Q�v�O�<�����.k$ϊ$�H��"&$>h6X��{�#�*8I��]�;U���J~�X)R�5�����MT�S!����>�ϗBrUn*�a<�}#�]e�o�tV� ��9>�A�I�I�M�_���&����8�C�q^J0�b�H��u�7���ʏ ~x��ʺ����h�U���y.�!t6g������91��Ƃf�Zx�����G�Pw��C�����l�5%G�I�D6�P�D��M��ո�{W4gj�%I����(e>��)��B|b��t�5������n����i����������4c�ً��=��V}rL#�*Ҿ�^����9Ó:bW�u��_e��H��{�����=�U�8����B��?6�=Tor�ԉD�O}�?�q���|#�k� �MtK�B��6��kV� ����M�c�o���Z���3`�^�]k�1��ipx1ְ"�� %�[NJ.'�L��k�Sx����B�+��{��$wfI[-�Iu	���2��-�	���a	����ΝoY��X�&B���{C5�j�ltG�[� ��hH��ܽc�;�k�H���dҔH�t�li�Q�y��}?:;������_0t�ϑDV�׳'YC��k�	W"I��ʏQ0�7�������#b�W�!���Y�x�C���>ⰿ�B���}��t��gn�I&�x��)ې��b�*Kt��k��{�+��s��G���,�&9�F%�PE���"��B����X�	�7����7kY;�H�f�ܚ�m�R_Ϯ��]����hcԝ�)�]Cʦ�!�a�_�a�߆��)���(r9x(��TJΈ����$Fզ;�3����]�A,N��4��|F�X��Wz����QG��R�]��{Q��5O��pX�
�)�]���;,RѬb�N��F]�Y�%��j�韀��z*�*3|����)�q!A���2��t{Hy�����-nx�[�^�D�*r¨(:�!��� }7,��C�b�>�#��' H�|��+b{��w}bb^�8k����Ѵt�t��*��e�񴣁�[�cp��"�84W�2�t���h]���!����2������[��Z`�a�3�*W�Mήxik~@d��3�|۫MCw�J�>�"@��#��W`T��>@���$�8
��-
	zJԙ�WH��9���,㟿��tp��8�ǅ�A�Ja ����#y�VcsK�#�헷u��ܓ��n����h�U�-�wWI7ӧ6e�?ݴ������;�����@ō>���x�,�`�;��vc͔%o������Z��m>��9}�%ǈiL
�:$����V���(EР�/+�g�s�5M����x?����\��s��|�^��u�l�h=4���&D�T�)D�kb��("�&`������G�*�X�S©�RBeX&�.)�]aޠ��,g0�N��-Ƥ���H�mBAN��ox���Ş��]w*��Hඪ����0Q�wy�r�6�n�J�.Q��@P�)Ќ�p�����|
�&��@D^�ety C��� ���ZV
M��!�=#X9��@�7����߽��ThQ�j���O*U=�mq!SY
6,� p^�,� IDP������WE6�jk�5����҆+NFк�K� (>�	�^�`�t��P�A�A��A����;�׭F|�3/4n>a�;_?��?R�z�T
6#Cǥ=�Z�l��z)L������m"�IA2�&�U �>�����.�fr�0��Pp`r�W�g�4?�f�b�J!h��2s��$�[ߙ7�Ӝ�dJx��h�$-�YFQ�K>|#&��/\F��a|����N���� �y�gQu�BC�$� �H��Zp~�*+}֍���iǍ�^x5�����(B*f(40e\秘�]����N��u��4јi߱�H�ϣ�%#�PG�䵪q��mTa2�;��[@�EBٚ�FX{�/`�Bsy}`�������yc��q����F](��e�\�Pky�7��iN5St�O=e��z�� �Lo�\�k�4���v����v���!��?�r�O�M���J;u��Y��&H�;����X��N��T�����RpYBQkC����"R�W��8��w��Y@��[�Q�Bi��2�Z�L�`���F������cML����V�"�܂x�7�*�DOIㅻjw��D$���|u���?R��6�$qe�NFN/)}�d��%�N.#F3�0g�{�[�S<��������݊��z&���`�L��mR�b����W�e��
��6ב��^��c�8:n[x�@=<$e����m#k�^�u���x3��cyo��Ĳ|��Y���2wB�-��*w(����"3b�cy��ӓ�$6O`9�A���M)�QE���Z<C�I�R�1n)�A��R�q���kt���*�D��B���
G�1��_pt�ٻv-j.�m��5�����R��V�]�y���~�������Q��%.y�JF�2+�^0�M�]mR�ٺv4c�c�Au ��
�}H��V��Ե�f2��z+H��	D�m��ώȥd�iޠ`�S@������a�?�ld�N��y@�:Dþ/�![��]u��H-�K�Ā����ٔ�hl�����Zj����X(��h��ůZ`�#���;�2��.Hc�6MT�b\:�����O���!�m{���e;uol��<,Q�aUN���Ut�<�!�6�o	c~QRz�5��u�����j΂~�]�88�c�bݩ:`OP��N�,7�Q�����B0����~i� Z��I�K��h���Zf}����h@�ypBG�\�NyK�DiY�XX6�>����,���n�>Df��,��������*X���߾���'l/���s-�4��.�[��f^��,�}S�̲k���j�p�#Μ��D�f�ONXhd���^����P�hg$��͍���x�����i��#���?���R,Xx�e����mS'v�gN5����v'j�ͦ��\�K$[\���)�4"��9���7����xf�5x ������� �_%�^KL�_�7������D�#�Ax1�;�-ic!��S����|��k��K8�⮞@:W�w���'�r���./�}
X����0u݂���H$R3y��\�5=�A�O1T�:~fĹ#;Z���ݣ�I���E��C��`͛׌H���M5����\�^�1�P$D�P}?j�Aj$òC Q����c����ő����v�6ӾB�&:�e|� 4S�����P���!�E����T�����A#k���+�9��ãt~���"�}\0 VA�r5�*$\��3�C���z3���Hr���Ղ럣wrߕ�k�?��>�넁aow�_=� f^�������}��a� a�)�ހmz&��� )��KG��#Do<��!�۾����(n�U7N�3s����=_$'g�<c��zJÿ"ۿ�����a�O��l�@��wvD�~�����_���RZ|��aD^T��������-��)�,���B��ĺ:DqK�u�]���CX���nj_�;���R(=�~
r�oXg�r������qF{��.#���86�[��Gv�t��*�0*��o��B���n@Qc]�v8e���)'�x�����\��w�"�5�<����G���*��>J���ل5���{�C�M#��'}x]!��?�z;ْ}@T ��o۔��;`��̈Է��.>Ǔ�Wg$OmBfi����ьf���){bCL��K�[�������3��p�dW2̭�H묋)1
n/*A��{Y�k�tj�9�����N�e�a߼7��&�X:���7*�������Jh>���-Q 7ճ�E%�� ��L��/Ƶ/�pg�0�$-�i
c��7�BN+�䡍-��K��X�%�ۗa̔J��/[l�%`�˾d���.Qk�V7�� �ȟf��
��~�Y��I��P��J4�v�~/�K���whm&����_������Bn��D��ي�ʃ�J��2U�܄I򶩼�C�ޕa%~���I�2��(�������@Ӂ�� �l�a�fR��ĴY�rqT~<@/|h\�N_�Hv���@<���w�Cģ�b� �~���Z��:p���6H<��1���n#^mG���U|�)R����W�<;�{�I�K���!�U��&��u6�'݁��]��U��hA@�
is^C�u|����0��h��ۻ�~�^�=}գ@��V˴yƢAB�������J��^�R�t�D-�	ЪO��o@ƛ���5}==�կl���5���k�8�<�OU�u�-������QU�-�`3�o|�~~�Z��F~�zb�V�s�h�"����F�j�Oh�P>�2{e��M�I���� ���<�Pq�k�5���"����nI�*O��]���"l��-ݟ'3�����q��ND�;N��w�Q���%E^�fC#���N.�
j,���8���KWM4�bnN��-9߻^�t��v4�>�����Me&�눓76�z��Ŝ��۞��:7[8㗙['Z�h�M<���[���o�t	�X�v�o��yê�kL������ԫ=~�ye6y�is"Q���m�$���]zK`�zg����	Xx�X̫����h)\ī3�ܶ�������J�%'Bx����vω��y|(~OաɠL݊h���Y^oDM.��Zw�'�7�^xG K��w�x�����2���)5c��Q���@�)��ik�2�'[R_�^�H��X�k3��V����5z����w�"A�:�c78$���ѫ��bGQ�7|̃Z��9~%ݼ��(������ �JC��M��jpQQZ�"�g#���:i�Z��o�dt��+�N!� Z�(ۜ�5����kQ+����Aw���ú� ��0*<�~z�����P4����a����c��4�������2n�j��gN�{���->Sq#��Z�[���=��ӷq'|����NT�6c�n�*�I�_C�T�y�3^�ý���1��ԋ���"�_,5��� w-O0�C�[������y/Ǘ�,�U�=�>Q器���<����&7l��=rP��â�������<�Q�װZJcӦ��
�6KXl�ݦF�?��Z�:v��"���C��E�"��ǂr�[��k�*�{�_w	��k�:B�P��DH,*N�
0XuHzx�(��e�����biN�^�N	j1&C�%� e'J����t�p`��9�R�ų�&$�x��5��V��v5)� |[c�w$Q���_i$;6��q�$~�g��2��*�Eѫ �!5	W ��l�J�Y���;>y�R�瀳5�(8�hT�&����+�W����5��E�C<�yC�P����繘-�旦��S��z
?��X�$r?������`�Rcp�Zٻ�M�^o�|��T��  #)�[�( ��������Ea����	� 4��M��d���<��}�e5���SՓ��N��g���a"�mo`�.��w��ُ�G�t�|C��V��=t�+OmQ�����͆��� C¾O�M��q��)�<�}!�_qF�Gc-�;<�;V*��w���H�üg�O����Y��G@&�R�4�l��oQm]_�?�6�/G����0n�Y�����r  m`;Ӥ��@lU�����2+��}���֠j�z����A.̱K:����E1ߴU!7�e�/�m`�12��V���������zZ�w��_��ܷ�֤)�8��ʱkٞ* �2��B�k�{��y�����(G�G!�BI�)����_)i*1��'�8�U}�b��_k���5�-y���,b>��r#��ۢ9��� �a|�s��H1�y�_@߰����׵���̕ɜ{]3RO~'��n���.�
��|^��L�;dqd؊x��Wż8�vZO>�M����}߻%��s�9�He_��2���q(�i��i7���)lJ�q�Hɷ 9K`�۝�c��|oT�݉��G��*qB�g}6�z�swE�Y��|P����e�E%��!'v����~�a�~P>|�>���w�Yv0�8�,��_]��W�����}=PƟ\հб�ߏ�`�����RL'�?��0�Ѯ��zC!Z�b�O�'#�a�rA6΍�/�<q�����a�I��1Q`���$�:v�ߞCoH'���K0��Eqb�/\1�A�����<��m��+����.w~�p)u���k8�U��5�"L!!���"�z��ʹ�,^,�#�,=�.�nbu�2{�����z�d�O^��"S�����@.dP.Ь�d!q���sEPZ�U�^�#>稤/u#�8�W�C<��b��r��ֿc܅P��sJ 2��[g0�<�:�i�:�����3#	G�"D�n��ﰣ&�W:�$q����5�2E�	�w+��7�����(K�6��h�����~, O��rw4��b��BdV=&�𳱰8'`�N(�J��j����2��l��f��r�u��E/��Ӕ]
�r��a�j�$���6�>$5�,QJ �d4t����&���ugg�#<���Ks&ե���XZE=S�h���e���ۥ�#�Ԏ���`�x��Pkeh�:������oȌ[]��E_����0�h6�k�|���׬b1 ��P�ϑ�p:��sU�_X� �
<1������m�n��;-x�Q����봝KB2U۳6;��Q� 4F�D�Z��� -[�	M�~�R;5���g�j�T�7"���ZV���K"��{(zP
����U����g���zW1��^��:�{m�+��H<,��08�͏V�~�m%�
Ī�AǾN%��<;#ulSP��Yg�}�<oR��M8%��߿��d|���FĿKϡՉ��0bY�1�wX�Q�*І�!������	�jQaw^B�x�� ʮ����	�3r,G�G�a��.�Zh���wr��qڅ���n���������Y�&��"H�ʱ.#��a�+�`R��i�k���
!ᴃ�I�b6��H[�ӗ5�ۙ����Mi�3-�^����>�u���lt�U1q��Ok'�QP�s�d!��K�	Uన[��Z�Oގ�YC'BL���գ��[��F4:wQlA_��������3.�	8a���X�r��U�Å��ʋ�%��D�N��m�|J��JPk
���q'�TM?z����cS#@�Y��W1��%5�U��X�"������7�g��aر̲����>��QI�pcR�o�a���`_Q9a�%*W���U�?����.����M ��+������KG{�»Bʏ�7f�}�U"�<_Ǻ��'�!��:�[���� �,�-���|%
$�����xm�6]I�d������Sڈ6S�>�e026��K욝��7rۋ��,�;����vr6�([wG:D�k`v�e�4P��a/���ihi��4i���bL=�»��Ш�#������̻Í����x2.M�!�6��e[]y{:�E�Tx5.�f�W�M��@�%�Ř���7n"��7Jny+�h���6����+�Y���IU��L��E���hW�B ���w��{��%�+ʏPp���т���29�1�/��I~G��5 ��o�+������?$a4��:Bh~�r���RJ١),'������Y��Tz�a#+�[-�iH��,�V�:�b��c��\[��Kˋ������ �;?�?��~?A,���O4�K��&f �»�D�2cݼHr��z�}a~�)E2B�?�U�e����(�h�8!o� �o�Mª�зX~(6҅M�4h��r��xxGBn��y~X	��\;��X��j�?V��k�����h�Q�T��Y�?U��"��m�$d��)i��:�ѩ��D�N$��ŉ�~�H?<�#'�Hd�� ޹I����擔�i�_o[G�s@�Lٕ*t"I�����syA�1)��R_�N����V�,��L<Gkh�+NU��@�Ϊ\
��e�\�����)���}W���DiR�aU���t���A�y��A��]G���E�3�&��F����*�|��1�R
)4iYA���h��89^�J�>\�3j6��@bS\��p��k	eV�p�h�&�m�J�уS��S�~©+r����qf�#y�nY���dZ�Y��S��xY�' J��6>"y���e��91�D�������\n����T��.8�܅"d2Io�����u6	}�	@���~s�[��P���0���PJ��V���nD!~t�HY9pY�Nz���  �:�jW`�):c|	0�ljE-x*�4R>=��-��A�(�x`�$�P(�7���R?�"����x��FaV[ ��9�P��$I����U�ɏ6A�Il�zVu;��y5���ťD܋�_i>���C��b��;�6�Ņ\M~���"|a�YTX��6~� 7�5ݞtW[�wx��CB��5%��S;$3>�؇)�nsl���d-��f꾨X�H���L2]����_���4�լ�l9�fh)���Z6��O�ġ��ZvR�f�ά����� %fke�����ha[���!ކ�ѱ�ˉ��v
�j4��4SZ�#�Ř���F9Ω��ȴoYX�Z+B�H��� h����@1�+o:ʃZ�Q�˻UP��C^1_)���۴K����!!�'-"�J_���|Z�ީy5���a�|�ՙv�'d"�[Y����ԙ�.�~��$�3�f���g���+Z�|=�|���+�Iu��"���X)�X7C��)�|�fN���2�n� �ƃ��,
	�WSLD�ݯ�\A��[�$o�R4�ł�D�oGv�lY���)�3�/a�'1.E�"�AU�!��C�mp��2��;O@�#*ê`�{����_���Y���,wl ݪ��<̛��oR6�S�;�$L��5�7CE��P{� ��d�(�n���x-�$�3��g�ʝF�>=��� ;��4T�e@�!ʢU-�C�鮊��\U�b[�ȋ�~��e�%n�`��rvo�Ը���syB� �.��a	&C+l��%�v�5�$.v� �C�-�w�O"����4��(7<��Z�?J��<Z�%����Am5w�fchk�ec�	^�f�Ǵ�8����Z��~���*m�QB�=R��Yy��6����݌{l4
T~MK%��*J����oD���-�۰�_���Y�Ak����L�a�	Һ�s���Ϗ<��hA�� 8�ӈ���dI�>�� Ղ~��l�$�pM���3�>GZl��܊6��(��Z�M����n���ב��#=
����R�Α]3hc�E��gV�¢�ɻ�-6���u���$�8��]���N傑ON�i���n^3B�>��~����"�A����e�&S�Լ��c�8F�y!�/�ZF�1�a$����gh��!K=1�hI�oܕ� &�w5���$/���A��]I��R�{T�zkx�V@?����	�rl0_P�5,����U����s�40��������?++/��3�$5S�A�����GC�[������ -<�e}�pUq�
Ϊ]�軚����_�xTzl��Gtp�E5r�n@iX������-e�Υz�떔��Rpr�Gv-�x���:	q�Ve�}Hv�Y�_�ك���c���Q�&���L5����!�� S��M�����Na��f�!�E�V�P�����Z���Xz����A���o���59&����Ȱ��1CI�7;���|����`/5tt��u�"�X�C���S�H:��F�B�ɑƓg3ޮu�}���D�f&)ܠb����\(��
�{s��#�u���Y�`{���'��yثŔۛ�7��I2	��c�&�ZB%�Ŷ�G�D��O��oJ>Jg��H���T L�=��.F�ΰ�p�~�:�NO:�9��d�<�5�w�� �/B��#��*CF8�������������:�r߉:Oxa�S64zO
P0"`k��yO׮���	�|��[0���{)�����쐉is���O�Vl w{�McK��������&��Ĉ [��	JΔa����b!����.�ـ���*zEt?ȭ�*���~&$�d%��Zh?^:��Ϟ���|���Dv��P�b��=%=̗C�nUQ�w��G��0�4H6o�F"|�̹��	O�DYlO��qfg��_UOv ��V2U�1/���v�<��=�F0A�r7��$�1���r5��O2Tqf�������qK�z��RPr�֦ÜZ��}�Y_�9%ђ
C��\I�/B�؅j�V` �G�Z5?�	ˮ}�)�q.U~a��/�����S�6Q|?��Z���g���6�]�=�QY*�4;��~Ҟ�c��0��O�m`L��S�ؖ~�'�͒�3���A�$J�rO�,�꣥�Gx�R�͵2�A��	�&�I�uyM�E�8���h���d	�����/S�2��8胍�J�u�:��k��;�y�nhVa�A�>ء���٣P���So&�f���o���g�5��o�څ})es���>���0�}0L�/�aj�&:�N��鬵~���k`�<�DKun�aX���k3�J:��ng�1��b���:���$iCſ�i0v}(�?\f3���U�X,�d�@�Tb� �.�vLNW��m �Y�n{r����J>	�}��Ć�����k����)�H߻�E��G19�B�@+L�f����vXx��Ąf��adn�����o]���t��0u�&&S##Oz�˾��nc����71�o�΢9���&�c3�V�,�,L����oY�!����(mɰ��,�h���7ˁ�߶{��oo���s쒿�5�v��(3p��G�@��ޢ��e~©��fά��,����Ӑ�����dcǜ�K�T1�O�t;\�(OO=9���
�m�w��v�g� �Q���:'4����(�	��;)��cH8`�z�ÛM:2X�X�>R�ÄW��@���X޴�e���,��=MvF�FÕ���.`�8�@w��o�(pa���,�����<3��o� #Hx�I�T�Q� ����߳֔ļMj��ZbV��ikf��{����yZ���F�h�w.ܼ�9Sm߿�H_�b���]���[=Ǯ
Y�)N���Gd���D�D�;=�y�P`����O)�T켘
�O�]�j���� .��07��������dAxV�J���Ͱ�x��ś������b��e��OJ
��pf|�-чP�	(����D��� T���Q�/&.7�F+��>�z�"�^�}���h� &��"��yi�?��~C����[�1�"e��ʘ<��w����b+Wn�L��{RrIH�V��<��C��xJ���|�I<�_�װ
��M�u�!WY��ȼY�!�)�W���}���R2��TR�$�VJ�Xʡ�*X4��j��z�\b�%S�V�c
Nlꕺ�a��O�lU<�rq�b��@[������>�7r��D���c�?O�ǔ���(�g@�G�M�cT�c�����b�lm���	���6�ƴ���l�M�Q�p���%��v�Xj;o����4Y�@�:4���3ք�Qn�ALO����O�4�yMua�T�Ұ">ov[t��![b�uHK�Ryd�;+gλw��2��0���D�&C��d^]�H��"Ԓ11����qi`F��a��-��[fB�6�љe�y�Xج8Y,�?���u]�e�Nn@��iݫ�m�B%��$]�V���|{��/e�}y��e�MV�$ ވt8����2�HN�x�f�cv�}K���r���Bkr�I�O*�
�*s�@ߡen����Q���N0�Gb���:0� h��#`�)��#�ɷ���9���*�;#���^�HgU�#W�lM���*�T��x-0���X�5��mt�3��'e(�g��O�C�],�7ֱ����k[����=&��.#C�8���M���Q��8X\��8)}�>)��}AσD%A.�.R�[����N.$�z@��3yf����iĭZ���&��l�ژ�7��<�A�@�火�i~�$�_	ϸ�ũh�RwbȖR�b�L�Q�e˅����8�:��<{�{/�>@�An��"w�<,��5	z�z��Z����̷Y0L�i禁}���oQ���rR~�c�������J��k�lCho��{�yn���b�ã���vt9���j}v��ta�f�6��?2$i�X���5D������P�%��W`M#�r���ڠ�Y��DG�=�1(5��.�P��=����4�jR"	>�MT��vA2�ʀ���ϐ�^C��^���T��k>�J��������ZL�t?�O����.��Hm�� �/��$#� �r,a\s�{��;���p���u�8Qbb��s�\�V�ƶ�&������\w,>�J��ũAz( ��p�j�֕8���ks墝�Q;j�aw�C� �S����SJ��`1�8��r� �zy沵���.Pw0�<$ν��U|�F�č���R�O��O���%Gc�#X�� 99��r�	5���\5�����F�f6�g����3�hx�ʺ��%@���7�%��u(aó���D����PGh[���}��7#��8և�a��o���5�>=G�!
���<C�y|�-N�1��0��FJ�ޚ���<i��~��	?8E�ƺ�
�۵7�o�5���oV��3�`�@�	�a�x�e)�U{g�5��x��]�<-����ʹ0|�����.,V�Q�в�iL���	�i�&p*V����s`G5H|��-�<u陑?��� :�!rO�A���2�<3%b���2Z#�QV�&����N��i\D�?�S�d1	�c�����D�͍-z��Wfk�����9�^Z^��D=�����}�Vu�Y_���evCn)�o�^�s	LQ,�2�"%���"k�_��ݾ��,�A�Rj�Av���H�ѿY���f?��v��gL�Lp���q�� ���s�nW��ij 
a���3E] }�į��j7oF���"��v-��r��xr�Fѧ���N�	~�塲�:��oQW`�<|�f�C��/c��_k�S���T����7�H>�H�:�)�p?)ыQx�4���N�(�L^��hp�P�������j���*�=�����r������+;�LǞm@]F#���=B��.�7^�`�"��O�љ&�_�^v싯J�O�Oo7$:XG�R�jBp�Nr���q�.n��@;s �,f ˺p�̫�N/���_Q�,�P�������Z�ZaI�
�T[���.d�8�91�ak�3V���I����{�e�r�;s&�!~#L�9f;O#�� r|;4Zy|����&�
<�D�m�j�NV���F�]Д�9�F����ڝ��:����*)��O�#,1�����o�1�u�������Yř�tg��ܨ�5�'��t6��x�F����g��}�@wxk�[�1�=�|�R�	���2�����]��K�%�pA쯊�dQ�� �<9�d�M�f��f�f��i�&�+�`�C�4Yth6]��8rP��5�B�!<�2i3�n�<pr��O�C�H��^3OC;W�c�,}`'�7�l[���q�Q<R��u�f˵�쳈��_d)C,�>�u�R���,c���V�xM_�n��� ˻Գd�Zz���=��D�ȡn�Q("ii��l �b�厜|c�*��T���&�'rCA�uy�#		�H��F��B��*���6%Ln�����Ǧ�w�j��f�yYy���궈0���q=qE7�9dܶ����VH�K�a�'s�U�h�OЦؾ}���\b�:z�|�S'�<��='+ߟY�ycsƣvZ����%�R	��Oݠuݪ���>��#Â�z�G_u��
���#�,�>h!�潯�u�c����g�i�qͤ�8/R��(�����W"�����裵k�Y�ߢ�4^����Js����8b/<:�"�,Hf�b��=W 0	��Z��v֤(a�r(�t2�p�x�v���ޟ�V���.����d�x��~F���X ���(){43���_�H"��s#[h�ʤ�Ƨ���v�{nH�U�7R����Xr�]��0?�q�d�Ȗ"���a��PW��;�kM�&���,��,�K��YLhuxS��X��O$*X��&�
�#U�ƒ
��y:�C�u�|V|�+���Pǚԟ&���Ha�Q#��U�����1�Ӵ g6�%^C�k�*�0���퐄�J��;_.�(��ۯ�Xd�T�_XM*�\�UdN�g�1o�M���S���>�I�E~aQn?61)��j�NvTF���'����ԫNgr]�]���>��S~���Z�|� .{���q4� ���ŝ���%�/[�� ،���^�!��U�	
���>���Hk��<z�2y��,�_����<�����*D�R�N����p���L���޿�0�H���;�~��\M����S��e^�����k��Le+å�1���|����,��+K�sW��l}-�R�e��ϢD:k	MY\�0��G�����ҙ/����W%�aj�i�lL6��,��{{�U�R�fA#�`�8�/щ��S�VJ��J얥�D(�T���dx�9qe��÷�F���7\�rx�s��Ӵ��1���k�+z����+*\�q��~Ȅ�;g�W��*�f;X��y!�tn� oh���s�����\��\�A�'����r']�PkC"��B�.�O���:����ē 3�k�}��,X�/ѴE6$��=��MW��w��6�+7ԕvb�T�+K9RK%��Ď���5-eT�}Qb��HY��x�h���.�EC�����O?GE{ʽ߃E�1��+Ė3=��`�*9m jbx/���.�4������a�:�@��	�[~V��­�[-��E���H���w:aK�+l�iK2���Zp1F��Q(A�H}BT��58�Hl(M-�2c�e3�0%7�����R)]�*�#u7��n4N��dm
�3�n��~5*��8�zD�C�Q�ms�����?��GD�$rv�B��J Sgg�e�1H��8��8(ʏ�:�΂:dظA�-6b1׫j�~i9~�����QS��Q<l��-�&~�����#�Wي��8Ҕ�Y�s���qȴ㱰�sA�z��;��nі�"E�p�X����Q��f��@.��F]�2�W�ҙQ�M;1A#�1�֭��K�-0:v*=�['�$��LZ�{�Z#����Ҝni�����U�߉X���欣5�ƽ:/���b����G=U�􁣑;�J�g^�iŃ�)+��;��>Oj��B;;�����j���例����H�MT�u���J�0>��E��Xf��Ƅ��)���
lȘ`*�dH���ۀ-Z���d�Oh��?��=���)t������w8ua�0����[Gي�u��x�4�@S�E��%��5 ����q�S�
&j�A���*��:�ť�J�z�^�:�;��q����t(�B�d ���>�1J�Y�`+���M�tv�����3ߗ���\CX���kcLK?o�G��u�5�Yᴗ���v`��U=�I�KOr��|��w���AT��S`�v7��)10�!c�`g-���6���1����[�D״�F�8R�O�eU���ǫ�ОyB���̖��K�8;��*tVav�N�h#�
"�e�J�������
�_��U춚������������uND��RRv�i�%(�c�c���7,�+Zc)�$�����{�s�i$���#��w%���wQǁ���3�A�m��<MK�{�I�K�F٤�c_�O��q�[�ԮF[0�9�:�EVH��j��� �yKb'OQ��~%�F̎T1��bR��}sr�E��Ut�I��h��YdZ_�&�nH{�+K�~����n�M��PMY��p�+�� ���ho9�S���m�4�gٙ��ݚ	��&{-k��"'He{pF��`%��]l�`��v�E�ww���0��/�3!�g:�hp畜���~HX*A��u�I�ƺ8pa�bf�!4�F>����zۢs��1��+��w��O6Q�N�͓��eqk�`�jTM�p��U/@7�+ԳR�GgE��)<���ap�M*��wk�~H ���2^k�%�Υ��i��gd��=��n�f�2F$
��:�pa2"�<2R��{힄;-�:s��ˤ�KJ	He@�c^'�A�G��F� �	2o

W��f!y��V�N4b��:�`ov�?:��u5N���N�J��ؑ8׳dd�����P�N"BR��iE����ia��lq��(7@<�k+�}�I�OA����QJ�Ė�R��(jIc(�!�H�9RI�8{g#�lH0�A�3b���0/��0W�!j�	�a08�A�Z�\H�O�d#7n����g)8���z��I����D���q�vt�ر���}�֊�s�R�5�����|0�B�$OZaA�@�X^ErI����zIm��������G�.Z�"v���~�W�K���V�� O���c|Z��p~uIiH/�&�D%��vE�	�ױ�(��W���x�6p��էӸ��e�jb9��CR���nrZˣ����e��>J\7��B�d%)�'ΰ[�{����'�s3�>�����$����L� m{�O��(b�TpM�5�7�fA	�����(�l�����FC|����UZ��k�;����R���U��j�t��>����x\��-7�pᣃ�#��V�\�Icu>��%�3��Z��m�ً���e�iPN x����y��`��=x�y��}�Vж��a�&86����T�au��0������~�_sB��V�7>�	g�1-r���[U"W����c��"M�OC�>>�����<��lY�}�8��]ٴ��<��ͣ���=�R4����Pgi�졛f��,�Ӭ��L��#�yI�R�u]`9�<R�5�*�*[�(|	
i%�QT~xQ�Y�1Gh���_�c>�=� ��[D-됮p��Y<Ą/ò������"*�x��v�?�|LD����<�6V���qp�<~|v؆̎��N(�9��FZҷ�ƽ��V��4�ѕ��zɦ���	�pG�=��9�Z )�3qX�%@w��neb|3��8�ڗ*���^��~e�@��XS�+Wo��|F#ɒb����T0�]��G�4�K�� ��]����W�MT�!~��[McF#o^����l��K��֟>P@S���W��e©���Ѵ�}�鑞%��e7�Y��`���1��mao�Q"
i�Y}P�w���9qx�l��[��b�\	zԦr\�l�����i��+�tEm-ܭP�BӔ{�����>�4�\����?&�=��	`��2�i
����|�x3O�c�p_KE����A�t��ꙜHE�XW���<�[:Iv9'E����2m����",P������@i�FK���%��U�QO�CIR�*ڲ�3��{�*��ӎQmV�@�$gXF49[��*d��
�8���"\M�ZP]�BJj��h*�R��^�W�dټaC�5?KJntCv������މR�#��^���Ğ�3�ע�f��������+�[�R���aQqىt�]x#�J�l���t9�OV�f����^�� >Oyhd$f���' �9��חn�1���z������K,U��!�����.ک���?I�󝴨<�1rEZډ�� �o���BuW�-��F�q��:��rzB/ߩ��'k�w6�5QHDm�#H*��,5��{�"Q��;;�DD�.��sm�\��c�^�Y�rd����l(��L>H*���H!�[��_I@��� �P�l��y�E�$�iҲǦT�ǚŔ-dIM+7���N�cd6j�6��3���\��6V� ))cÊ(�p�sa�#ĂL���̶��AS\5�t@�تK�@�(\/)�8i�����+���x�3UJ:�/$WP�( ^�b�ʼ�w�#��a�������E�P:E��_c����x���6�2�T�m�}&����(���ҤC��`�y��C#:k���[P���%���eI�Sh`6�a��c�v��L�|�A�<��M�b�1[c�MΜ��&��1���μk6�&`߬��t)���*���v��(�-����x#�?a�@�,^;%��3c�Cl�8}&��cT�r<�r�{?��Xb�5�4w�q7�̧l���!i3&������w���Wzov|����s3@��(��3_�j�u��!B�ԤH�W�f4�3u!]L��A���0'�I`]��6#F�w�h��p�`���?�D�}ݺz?�,"`ĳ���;Щ�H �y����wO����sl2���»��g:����o��ؕ&�<��rq��C���_Zo��!"u���$��i^ڹ�.�8��T�ô^���rV�BL��п���]F@Л0q�\l�m��%W�'$Թi�}Af*)�RF���ҭy�vhC��So"FBHjvшyo�� i>6��Ƒ>NCH�1EJ�����NS��Ň���%��w��uCKy�1��hNѵ��[�+��㷦$�s3�A���.P��`R��k���D��:�07�C?d8)��!o����w:^c��	�A�B��?�nL>k]�=Ft���Or➻��N1�:uƼNv)���H:wb��~��O�!�'�~��T����z��05�0��,�F^�cW,�6q,�-q0�QX������!w�n08j�����8��`�.
�w����T�W_���)�z��}>�x��|�Qz}��)���K>}�h��5ђ%.�l����L�E�:V9��D}�q_Y�Z�:�Wx2U��[���]��_�Ӫ ��`fǄ�� �dafK���k⻨�?O����j$oދuꊇ�mfΩ
��7Մ��k�ޠ��Z�c��\v��p���@��l2Q�c�b癞V��3�m���U��w�C��PGG�-�,��%��J�Ĵ6b.�f(����un��7>Qo.�:F)*C���c1Hz��3��`�S���h�u<Ç�ԜF���-�j��x�f��|�Q+m��;)�����)�F�*8.h{M��*J$�ME��	�s4�F��m$$�%R).����a��M@-�_ �G���0ѯ� ��М���"���3�~ĝC/f2�R՚��uW�h��+�jJ~��� gP;hWpT�@�����hL'~J)��|�Vu��FE��AK�P���	v���m���щ
�Jh�9C���)IC���K��l��=�/��V�yH�F��S��'��8��%~�Zo��A@���\��7����Z���؈]��A�zeH��m��%���_�&���&!��P�W��9��!��h�94����͓����ם�7��"<-��ݰ�m+�?��1�
�>,�K� �Ő9@)7?wݪC�
tl�f2���KfpjD(�k��+�� O�nVY}��):��\E���aA�Ma&�	M@w,�_W�g�ћ�3(3�ǣ��y���i�Xv4���$|��	��%\ؗ
���0�F6���χ���,����A[ҟ��Uq##�&#�V��*�q���E[.��j�\'�<7�6ψ¬���:afc�.�)а���I4�]�̥Іj�9�/}�:�(I�����6up�$.8D0�!C qCy �����d�k�s+W/�1��U�l�&V�A�򠠑<���/��(}i�PP�0��_�I[�l�߲E{򟨺��N �7�H��lR���e�=�UT|�0MTY��	��\�=Go���D��7lZť�.)th�~�`�z�\g��v�1�]��������!s���<�Ep��}>���8J5W_�5�	�{C��#.-���X]V<��o�\��LNډ����bh=�np���*\��Y��*t�oH�/����PJ�\�cl�5G���p]s�++�[�]��)���r17J��Ԗ�a��WR����V���o�ۭ���S�t���
�"-��)*�
��vx�S6c�4�H��!�eS�E�@�s*W�N��X��b�UJ;&R'�q�3�����;XU�U~���F��st��
p��w�V���t^����+�	"�����@�U7�)*����Itx����ӄ?�SҖv���8Q�9ˎ��x�_=|w&�'@e:X>b:�}�k&��<�^�u/���jR�t��P������(��r�\�輆�U<�	��M��&0���G7SU(����aYI�S@�>����M�m���4L0�� �kK? �h�`�GxQ�f�j-<)�R��G��?E�f���J��|)-�De!�=�����>43��E�� �$�q(��a��ޘs�M�R�2�F.�N��"8��k��b������m�˷���V�p��Y�&�K�~AƊq�"J���U���ƛީ���	�����9�˶�f�c���e{|�8�^���i�pN�'�o��V}�v�e��S*��Y��鲦v{�!�/�c�W��tDb���M�aP ���S�Ng�"H�P�1�Gj7�1���r�Ӈ#��C�EYJLy	
���M�vy�8�s֗�pw��ë��������rh�-Ԫޛ%'��ZA<h
�i�r;C��fnʉ|Nr��H���~�`�e[�Y��s�|�[��`��Y?��-�+����X�
�!Y	���z%�3���MX���Q�龧W$<;fJ����1u����b��}m�}:�U[$����ʷ��c��L�fA�5�q�>�N�-8 �s��PD#8
�;�N�$fCn�:2�_���1���V�ctF�`]�N3��6����e���M�Ԫ'���'�.7�!T�Aݯc�G�1�j��?���b�! ��qi�ŝ����Q�?�X7���(�?N<JH�vA�oq~k�˫�>�,D��o+�g z'��,D�j���g"M��[Փ�zSp�{C�D^/:]�;��Ղ����j)]��䍩=��E$�X:&"�ŗD��W9K,�:1=�(��`�7q��Ă�5\�?Y�.��v�R�����3B��e�Ó(�b��g>>�xT�Ie��ySΌ��7%&�AӴ����[���&�ho������Hұɡ���������o')8�&+�6�D�S:�^� Ԗiɂ�J��ϡ��%&T�&Z�"���v���'�(߰�`��#���jFo��b�^ڠ�^7�ٛfN��\�$���-��|�p'�@T���n�˷��T��0�R"��r�]�Um!wo�J�f��8zZ����9�/C���y�a Qܻ8R�#�{�~�š��h/�W�LM�j{�kw+��W���]~HC��
a�<��'΢�����Y>N��j��O��>���.%gz�]���]L��JӤa*��+�9����xp娆Y��ڧ�an  �_mǷ]k���Fj�wZ��6�=�����l��;�X��)9�~Ot?ʈ�l��!-<H7��s��D�����a^	��5F���2�ڐ��$������J�!o����O}�+��쑢o�|��r}��\�k3� ���9��rM4��}qÑ�FL�!�)Z�e��_4V�͊B�;�r'X���l���沤��L)�a����w�ŏSWSJ�f~�冞�l�֐�zN2�Ȱ,�)7���4[d}Iu��O!pABb��#��L�����[`�]N�{єq+�L?�nT�FL���$.�#
��^�/���m̰�u���z�<����z����LY�� �򕉽fY����b����1���6R>�;�kY�o�y|�.���ZǦ�.�P��=�q�3�9\��	)ujg�L�S���aZ7�#Ӈ���Moj�g�p��[}OURb۷F�� }�҈1��c`���p&�}��:��L�Z��ቾ����F��HL�Y���r����L��9,ѩ����"����q��Z��B�o��+b�x�v^��A�E��Ak�A��v���i[�#�����G����r���P��%�,�k��� ׽���q�;�֚���8���t�tF�\��_ԭ��E��*F�rf_��>�M�^�(/�p���b�VT��Cم�]&@��~�`��R{<#�c[)�Z�+���7/�9�N8������-���0�n<л�:Z
��Dж�����\���AVE� q���f����,��M%�KR����T�'�aܙ����L�c����fbU,>�S����8��]����PM*f�K�=��Z��pW����3~E��:5����`0ӳe��Yd���*u�A{z�ӫ2៊��kD�<�rI�!L:-��s���$HF��/eX��b�����p`�u���E:�O�f����P ��T��Pޫ�ќ߀�y��)HUo�GhgJ�@�NS��5VB`^R���.4p@2��Y�H�G�I�f����<G�/k$�0o!������<������R�p�L�YD��O�b�,*j�ĒF��y�֚�8el��7�$����9:�~�1��G���%��767�]d(u�>�!2:� ��o����m������1fA`����C��}{�[���fl��~%W�at}P�0��n�����G��S�+a�5�<���E=6�=>1*<�Ӱ���5�n���j��q���F(����^��4Y�E"�0�4��
+vcY=�^%J���B��:&��A: �����I����>y^�xV����pSU0�OQ�;?�&��(|�x��,4�(M��+Y�v��ɒ��^wt��,�U��^QE�?zv��;���3�REVcA��7Y;��MG�kJ�~�b s��ஔ��b��me��?��賶l��=��`����8l�e)Zlg��J2uy���������z��ӝsai!ؼ�:X"�{ �Gs��<����ʦ��S]ؚ���t/�m�o.��~skao.�e�H�j �����/�� ���tV���YM^�$�_��ꊭ7��K�#}G?�V�%?V���@9���{�#k�O�9`��1ee)���\du^�s�NLsİ��U`����l�S]P�U��bkP��͊Q�ꡣßvm�c���M��3yS�>�<����-�؜ޖ��n� ��V��c@(>�4�����j���c���a]�_ۄ/}�}52.��pl u�a�e1)�䷠G�g�#FH5�F4%�B��C�zXZ1d��.�ʮ�Y��=�Ϭ��'�V#Jo��ԶQݔܯ�R��'�<FU\��c=�D�3��|7��U�kA~Ȯ�X�}�߷V�2dY:)�wo	���HM�fn�e�8q�N6 ��K�[�.X���2�5-���_9s�ہ��PFMxE��x/��Yu��p^p����qqi%}�i�_���?���8~f��9�h����έ����%��Nur6�L������ʧ����_��������	�7��q��I��&�@�Yxn�z�1����$��X*ɫfŴ:���y-$"vXr�b���j	r� �i���W�^�8��^Șs�*��լ2ZX>�o�����"��jr��G�̳���E���H�Ip���R���Z��6��@�0���,�шQ�:�Pܴ@�)G��Z*W����yHCm58��pK�w�A� |���V��ЁRb��yi�C�y;F�~�3;�Jk<;c�"�lڀfwζ�dXq�
g
7EIU P�݂z8���$�kR쒗���52}�q��P�[����8�.��n�J6�I�m>h�e��ڽ4JJ ��c��+����F�k�;��T���"����̗�(�m|e��Q�Kl�E�jy�r�}$2;���'���w�20���i������������8[K�w�6��bM�����y��g(����$t�ɣ	�7��H��q�u���Ç���in�z�����l���� �a.	퉬��(S����}E������*4c�����5A�,�c�UE��^ȤWD� �i�q�[��?��s59nXGt�`�&P��^z��������-�*���~JJV�X����z��z�k�g��&< m��`��)P+j���ȷǶE��`�|���K2^W�`�=���5����	�� ���1L|��^u�?���o�gY�}%�od�~@bu�h욌�Sk�Ȣ��4�F��
�	
�I�F���w&���t݌��:���%&ޭ��u�9�XԂ'.�_�1>i��,�۞��񥓭�[��ȱ��v��hN{)�!�C���o�CvU��mu_�z��?��$
�׺l�4�;��)�򡞣�js+�bv�O�n^�)�g{�E���Rl��I}�)le`��"����/�~�~���[%�n��MC�!)�?����bV��{���%�*�Y�lP�V��K�i)r���~Z*�#����}��򍭣5�J�ٹӔ#R�΍�����ى\?�\��MnRè�$hۀ��*�.,b��	�������xy���������$9����˺�K�qO�T9oz����F&��Q����N��|�	�4�e*�҅uIsNIsqm]��~ތ��Ƿ�7Nh8r���D�.d�2�����ImQ�ʩ�&P�衭0<����4���SE����j�;T(7ߡ-9]+�>e �(�?��^����\���(�l�߮A�
��>�%U����4��s������&ހ���/�a%�;c4�v����-U��y�a��>��� ��m�19k~:����0/���As��L=,��fFy6�{��[�,��&��m�Ai��Oa8�Q�%6�>�A�h~>3�e�t��\;��2����M�Gl���푚���l���O��vLl��l���{���j���4-j�@��޵^��cg}��:� ����d�9ĥ�찇��ί|���W�7"���o�_5'�$�]�n����=�zF����JN���{ʶ�=.P]��T��@;�or=�����Nb �^!~�\ƭݗa�,�f��[��9C�}��˙�ٱykC0�8��h��6�o�V��b^ ��C����a��Zk��`,
4��7��E�ኛ�=$���T�8����@���xJXG�XKp9�S�o���"�ݪ>��;�D�i�G�����K�(�E���i���5�x4O�u��e�2<O��0�^X�Q�`G�	����"9,]%HWy��q۴+:�b�U=d5}���`�{{V΄!?���G�}v|4ۏ͆cC��X��x�4i4����^A�=ѩxyb��R�4�c=NQ�L�摪�#��<����-���l�M�x�/�\�tV)�l�o�
���L4-����z&�m߫�M*'W��*�Ќ��z��a(�ԣS�E�������		��|�Ks�>��4�s���7�X9��r�b���J*�zE:����%�������{��6���N6�����5H��2]�}�����S����_?��?�t�������@����9�0NE(�ҳ�>lt\Y3 G.cg�]�}S��X�A��H+��RY7�,��������5�3�*��%�wY�߲J�!>��sY�����Ia� �͝kN�z�p��9�Ƃ�z�n�N�5ޡErvmX@ʱ�sfط�^�iX��s���J��u
K��{�nX����^j]��l�^�`,(B,�M��0�V�k%v�ڰ��.bf�4-mpjk��z�<��/V�E4��RwQ�h����Ɓ�`+f�W�B'��]���~OB���^��̏�M#x�(�d:�����N6��r�^}��
ǒ2؀h���������U�*�䯵7�\�#;�G,����d��<����[C�ޭ�M=d:)D���i��8�y�_s���}ۘ�l��YU�8�zox�(āIb��m?u�H���Y\�X1���'����`���}�T`�_N����?��`�W^�y�AR�����^:�����D.���7o(�S/'	���N��Ҥ:��a��u��ūW�.h�r$�#�t�g�|x����N�U�,h�Z�7Us��wA���tL��cS>A�}w��#!(�����.|�I��:@�[;�C� �e'p��P1A��J���H+;ݙ������Xzݬ��Cu1A�����f8�KPT|�hn�"��ۨ�u�h����̓��o1NC���	#��-���"#�����+L��rs͊y�2^���j�{o�[N|٧{'@{�)���U��%����?��J�S0��L,@ڢ��"˺S^�EǼ��b����� x��i��a-�E�aA�<*���҈��WN���*��.f�x�zk�C�b�����Ćwʃ��<�V�V#"���,ԅԜ�#MF�?ٛj�>�U^��?~W��&&ʱ{��_d#�4Y�{c���L'��ـJ�'�����?=�`8�b�Dm����C�ϦuѰ��_�:����͎�,[��u�8)�&�L��T[4Z�8����r	Ö�l2[��ѱ�c;ԛ�
٧=�?W���?��4�v-�i�g�
1�>k���~K�&&��R�� n�L��w�`ш�0���Bʼ��E9��^�;Bgd�Pݿ��b�e�f�\�r�j;�!����
J�,��غ�j�cO���m- ����ƹ���U5g��_���\��_h�ԅ��)��{���t��g/4$��1A���¡�L��x����e(�-~���TM��A���ߡzw�d����~��-���;=?��&���E�n�(R>�^RJ=�ٮ���.$H7�����?Y��ZP �Z����K�E�6��z�C�h�J�Z=�doig<"��}��W:˒W�Q�pΡ�f}]�RF�Y�P:"���.���#�-���-����_2�
�K��Lm��ߴN����!���{�����X�E٧&���iêՏp��d�OE��mW���Hc��WZ������;(�(�O������|���>���Y"��ba�ō����^4��� �� �YB'��Y��$2%���փ��H#����[�i�e3�( �����`W�2pU�#�1 {u�~����{ ���q�{�^�7R;KK2����%�\�:�'�%妀�H��W$�YP�/�M�5E��c+�x]��h�5Q���\7���g��~�cK+aFQ��=������ѐ�ļHGSVh7Kes���6���C�R��~:B
xsX��=c� ����� ����%��k����#pd�E� :���]��J�mti�2��AF�bx���P1��q �a�6}l�I(J\v�b�X�����14[̰B%�Ho1��[ [��.7�e��4E;mz��ww�ݼ)h�9���Ԡ��`zI��e� �a�8az��?��i��k�C���~	����C���]�6L^������nO [���K %�7!ӝa���b�n��?�n����Ko�Ҫ��\��M-����ɠ���eۈ����9�]�m�rh���wx�W�_򈭴��ns|�v\WB-X�WY_�Ɣc��QÉ��?�,T_"�,v^������tYJ�Yy�����ajUz�#4��D�����@މ�S����k�J�[)�<�\�̝�KHSG�$[��t��Z�M��Yީ��~��#*�cd��:���1����䀹� =˪��޸���9h�	�e~i�UH���0ȢV4���S)��%���ϱ���sꁎ�[m�/f_��`�$"�ƺ�fg(��p�P;*��܃�P�[�������H�������L�3ʌ��'�y����.���&��~�q��+���Ӱ���2�9\��S�����+���?A>�|�k�P��C�Q�7�����m�~���]�Z�`���0�t
}��@g1殮�Ws���Q�RY�e����d�:����x����I�!	�b�{��F�{9eJG$�������g�|�����Yۭ��S�RV3�I�DD����Mp�h�S}�Ӂ�tx�����������:��C�.��y���w	BEg\�!a���oa\��/=�B����%v��!������gX�E�fQ
&���AE��hL��>��3ڼXQf������U�d�~[U/��RB��'e��mA �����E�G*�f|�٭�ۖ(����_>����ri.:x_nL�x��~6qF���c�RN�n  ��5���B���؅��R�]�e������Y�f�}&��3�:��-?j����M����n����#M�=Rӵ9ȝ!1��)?����\$}�Qt��;ض�)1M�SAS� �u�{|p�A��bT�w�f�L�2\S(� :�v6�\��2h3?�y�8����"���G=��̾)&�"0k�$���;�����J�����P��+�^,+(����#��:��&�u��-��q�3�=a')�nA�����X5&��˂��J��?4��2'ßT�Á�����GZyo�:D@~������o5�F?_�5B��:<����)���H��+裴�m[�hv��ujG�7D�Ę�	���Eh��Y>.��6���t\�d�ϊl�����)� �E�]>Uk�^<���BĲ}��7��Q��V�GHyR�aj��Ԍp+��Z��fR	�	�c�����`gA�qU�l��h���"����:�d�W �����~��T�ԝ�.�^&�^~�i����}�a��s�IFYwزn���8�C�l�W좘�?);�|�+s!�0��*��d�����c+�7�����=����=�i^���O1����Q�w%�Z����&���6���;[.z ���w;�5;js�:�i*6"E�o|�`wAy��z6-�����mu�����p/`�O�)��In�ߜ��'�D�f�AyF���o\Z�"L}b�S�k�r���3i�v*�.쵘,;�]B��vK%FJ+:r��"�L�ֺ��V��<>�P�˱a��ﱱre��^��!o���A�0�޺�����w=�K����c/�^��޾Qg-����@�I��S�iӕ(��ʚ�?.��ߌ�S�z)7^�V�ԃEkc���L)L�����z8K�I�ԅ��픵)�óh�|E��_�����'�|����A�vV�{�r�-Z	Q��~v�=�����(�pg;Qdn� 8��T�pG����G3����iZ\T���b��!˰���5:���+'�V"��Ve�$Lw|����еH�c���<�5|��l�{>���x��Z��ZQ}
6�31(CC�υ��}Wok�����˼O�y �;^���,ũ��~�v*�=p `P�q�
P��J�Lt�"�ϻ��.��OֳFu���=��[�F�����ͨ�'0�Hrئ}Hs� ���'�R����؈�e�ޱ�<�Ơ���~��^��q��3 �,�KP'�9O�`�i�E%�A29�`� �h�+X8��חr�j�Z�W:زau�@˪�Q֭`�~Y��;^�T�>���(�$�&����,�KL}E4�8;G�6���`�l\4���
ˀ.F�O$��3M����`e����n�)ۇ�+��Qv�gᕮD}n���Jx ������0a���1��tS!� Q`��j�Uc�s��C6��c24���٥Mb�lfU���^��Aw���0L{\/�:��A���>t��L�����QFLȔ�N7�.f����˦z�Dd�H�G�=�W�#��k�"�5��(�a���,��XTb��߼h��V��$ήUKzAuF�@Ә�*�|�&f
;�����rog��=Lj*�q���;`��~�f4�ޢ�o���|���\	�(q߬�o���a࿦�]U�c�1GM�G �̞�^��&��xy��HyFs���>~����=Z���`����v(��G�%H����_i[]��6.��r���`�=-�I&R�������(�.���뎴�{ڣ�xur�BHGu�@H�Yz�l\}�/�ƾh;��So�㲶�7��!}��6�XwH�����T�X���'�!�`�����
�>������+�؝�H�8�*e7X����!SSo��1����j��
�@"�k�U��*�"�;�=�`/�R�rx����P8�%��Cbh
`*��X6\����!i�}ؘ�F'���ڹo�R?6a�זeɐ?v����7�c�\��:I���c�����7ţ6�4JR~��>��@��u;�r%k��Vvw��(���?�0FsT��Ss;�{;�.a`�������(1P�:��N�m=�"�ų����?��i�W�Ь��П��Qp��p�)Y-��e����ö�� �\!�Ɇߧ+8�kN���8_U�Q�]��[ա�Y���`�٧?RKM��gHf�F
��jgJ_��m����Ip��� uB[��'v�QX�Y�s����D.�˛�5!/Â}�aE��# e�?�� 8z �`�7hgpLnh)�ⰗѰD���H��	�c�IF,�#(�-�5�����3�1g�u���nm�a�#�ȤN�Sx����'�4����zw��2��j�L�ɸ�W/�C��^J;;C��[��/fEv��D�;����~W�C�1%N�W���ڲ����*l����\�ɍ�iv���l*GuiZ.�9��eY-�o�XsR&g�n{|3��O|���n{�t��e�Kg+%;���5�d~�/ȮI�O9� ��u�t/�%7�M̍��K�f&��'���؟�J�{�$H
��I7,Ko��y���d�z���wx��WVK��`ẐbH�f�׻|?���nd�D!P'�wu��f��J�xϦ��Bz�r�l�:	K�l���r��ޱ4�-��o���K]� J4�Ox�.��]}>�7BN���A��tI������Kd.�&���#e�痗X�yb�vB%��W�$<�j :t���Q�^>eE{��(����W=A0ϡ(�L�������j��:0��3��2�Bp
V��_s���g*�����������ۇ�;|��:M��31�Tд��W�XO[�&_͕Rt�Ll�v$Ŏ�0Δ-˯S�S�_˹�5�̊Θ[��My�_\���E��ˏ�V!!F�e��8�^g���<
��(�A��N??L��0*[/��������Y�}2.�c Y�i�JBCE�Cn�w&,[�Ph,Q�,(�$w��y��1XL��K�W���>�D�-ZZ�!<���*ޠ�z�D=�2]�N��o�q�Z�m��N�����U�A�k�Hx�a*����8��� �x�kٗoċ���n��ף��eI`5������vx*SWJ�A({A?X�\��|�/�j��LV8F7�3jJ�	9�zy��m`Q�ğM=q2׀�Fo���GWC#�3G����}�m�� �?m����;��x;��B4��8V�.������ f���Z^aGp�{��_0uf�!���l���$:����4�a�Ë�.z9�q*�
�j�UP��c���&�BJ�����_��W�oȇ��Y���̭�����+J��8Y��m�7Š�1�@EcmV��v�7�!�u{��o�Ay�E[^�5JH���c\���ˑ�إ��2X'؎��(���v�U�8�ԯ=���=!;Y�u,�cx/��|����b ޏI&�R��,��i8è� ��ǝ�M^��pU��?m&�u�	�Ϋ@�����e���1��c�;+�C���ۮEޱ->}'�� 'F"T�$�h}����y���]�K��D���P��(-��ʝA^�6$��$���ߎ�)��L����J��҈���d.0����G��8�U�l�z�z��vbV/�
��/��/=�Y�2*{/�^p��?レ,@�}���z$�>�	�:g��;��t9�b�[D����{��a�܍6ؠK��S��h�V/�K�!qhF�~">�B�6��fU9�'!V�I`����\���U�����Zk]�!�����dxp��3y�ю�lD� �X �C�gF3�o���T����c�
4(H��{�e��}q�*E�<��x;��s�W/7��C(�_���bF��;�ެ�Қ/�~;��\̥����=�r8J��N��n�yc&�=�֘B�$�HB=f��L��$���:�")3�k��+�L�9��$�c���HZ����d� P�^0���\_���j��G����Z�m�8�}�
�v�������߇2����5���+DQ�B�* ~�\�d������\[8�\��3��w�t?H�� t�@WX̰�?�k�=b[hF��%�tVt�ww��llH-wO�'Ȋз������}Y]M���{l�n:��C3eJ�!�W'��]9~˵t�>9�.�, �
GI��g�����_D�$���>�&�'z'햗ݧ��[-��A��Zj�~����؍��$.�Ua�{�Y3Iv�c���"�(�Yn���{i��	3�\Sy�RU���vG2ۗV���J �o�ȅ�Qf�v	t��v�w��t�_̀�##K�i�p���8�ôVR�f�aɇ�$j��BO�V���~Ca�F'V�5]����2{�qڣd^��CI���2�{0�W͌�n��Y�����kОZ�s�4$�wDDU�\���.��}G����p�R |�F��_�D뒱��S]q_8;@�\�������d�n'U�?y��`���V������h>�y�;B�	��Bh�	;K��Q�#5�n������T36�2����Vf�x�6�O�F]�Ao�.o��i�K�'M���nʥV���:`R����S�WUB/`n�� �e]Q�/^V<�A�oDjҴg������������ ��۵��ߗk8�w��*~���k��Y�'�H���ڤ].5,�v�BY�].��@�3?�G�WЦ�\�y����L�����&�m�߈�"���-Ze_��)�۪�Az��$�g���S�ܢm��<��mR%ROP��{W+��Lю��|C��U�~�4
�C��R�ԩ���Nq.�����2b&�^4 ԥ>ʜ#m/ᱪ!{�w�9h,��hiYo�z!��*��Xڜ
]��K��\Kd�їg�Owy�$_��$�1��iI1�Nv���$�&�w��p�=�u5ԉjH�uЁAF#����o>�5��)b66�x11���*����L�W��]!�P/BĆ��O�W,�*�Z��QaĖf���k쫶n���S&ת\�9eǅU�r3u?�BJ���f��r򥟮�~Q�ON�7wr�����c��I�<I"���-y�(f>"��O����,'o�)��Z������NM��|�$��x �.�E�܈upW&Ƒ�f��%(�,�ak�(%[S�{'M�{//6��a��zX����1t9yRm�{~���w��B�'{���x��eyj�䐵��s�ʾ���?�Y���/� �=���Y_��q1����/l'����/f���u:s� �I�S�e��HFȻ'1<�,uh�^jO~Z��L̚a/�����qc#j���8���hڡ(=cWF9>���
�2��P��_=���û��X�������-��x�̥�_�%y/�����Bj��,�R�������&W�S��WYƹ�>�b�ڴ�f�"�=$�D����(E㙌�Of�>���kP�1/�lY��1?;𕇭֗8c�d�aϲz�$xV}/�xK8�9c-��]�&h��ES=+Ι;�!�*�{O:k�r-�"Ni����u�h��[=��2�@9�������4��J+{��ɐ����N��1_��&eM���1�n�3�PM�<���ܦv�/R*{���9|�u��+����K�foZCߵ��0#�g�7��t���`mt|�X+*S&k�C�A�iE�!8�!PPq��Sr��T*+�Bu!>��^ȌH����,�"vx�-����@'��3�h?^�'c����c�`��@��S4�	nc�8�J~�����D���(�'���
��LJ¢[�f�wHN�jzx2�F1��1�Q0���F��Q:}%n��7	����p���m"�q%��6O/�H�(4)�HD�1�5� c�븱iT1���B?��o���԰T0]�v����s'��*#ɻ�ء�i�o���:�g�5_�Uu����T2Ӝέ���'��E@��)��c�{U��Q$��}�.a��@��" �XTa��/3R��-�g��ʇ[܏�>��>]�p�S/^���H��aLܳH�2��9���"�r��݃'v�����q�,�B�h{�t WO�g�U��O'2�|�5f������,q3��Q3��_4�6�RF�#��-�Љ�}�EO_ڱ��p��+VC�:�8��p�;��!�E(NB�F���S�YJϺ͇�Co����V�8���BrǪ�̅\��bx��t�y�,�[����>�0�?:on�ږ���U!Z	N�솆(����P%p���DC�>*+�f������.�p��?�[�d
uw�5�M*�K&�m�1�(tי]�J��UG}�f-�m�Q���=}���U���N�!��8��Uj)~��.u�©�̢��zn����^jx:�(�\Λȵx ���K����I��K�7�G_69!�w��?�q�& Qҋg	Y*��R�.o?0~��R�:Ӿ���9��'Ig_PEǲ�L9[�<��_��~A����`}���ܠ��H��'tYP_pD-~0�=����U�����U��咺��g��R�6%����F��w�[TK�.�<�]e�yW���^Հ)4�e!t��-��A���7��ݸ�J8o�Rv0&X
t��Z�S��L�O�{ ,��~�Φ40�у�̘K�"���+�w�|��H������BNe�&�56���
n%Z �B��#��T��!�F�r.JT���}_�i���0hN�2��T�� �@����b��Xr����$5E����[���� dv�Eյ�r�m�5��5���.��j?���ݛO�Ȧ�L��c��oY P���0H�z#��Y�Z)##����g�:Z;X�J-9�T���|h���Ȏ��m����Mu�4��1��'u��`��ʚ" �ٜ��-xp3�ɚG'w����7;
٠t�4����#j���)������Ib�����5Q��x�mI<e�;]	8�b���\�}I�.i3>���u�M��D���t��?%B泼˝5�Gp�e��u�F��$��ϐ����=� �#�B(�P��2f�`��,��T��(�ۤ���4�ar����+d%�|�i�f�xw���k���ëx�N@�6b�ò�S+t~/=��ZS�)$�ⓝ5;r>�j��2_�HOf@��P4^N�F݈ ��DH��I��<F���G��} ����ɹ���*G4|�X����	�e��N5{��[>ԋ���Ҳ�F�0b���:{
Y����b6_�Y����Ȧ5qٜ�X�,�s.֪:T֚���B��Ø�����:�w���2>�n}N A��W�}��$�~�Z���j���t���6�B���%Q��?��;�L�j������?��o$?�PA
XVϺ���]�O�YwH�AgQ7"����~�ͺ�_�A ط6X��<���?�~��0Łv�К������W����Ueѕl�O} �郤�m��
�)���)#���s��\��$�,����ѝE!Rw��
��(��gH��h*!�tX�:#���'�%S�čC84��cI?�u]w��s��R��8�h��b�cL%��/�\�A���d����&���K6��m �μ��F<�eػ��u>�+���d�YI�Kl/-��e(��o'����Ȗ��:�+��,����+��5�K���c�I�=��=�>��Wi4M�Z�4�QX���\�� ����b�Y1�A7%�%��P��mO	m���?��T��-J�	�6gY�y��U�>"꒍�e��$�RL@�΁2���s���F��dͤ4]�Hiߧ'��hn�013H!U�e����O���s��|]%�ǆa�.	X.eK���p�N�s7���H��Bg��=n���%aj9�R�	��jtF$�1�Ω��I�/6�	��?�8� v�9[����e!��m�����oԟ�py�_��p{��"Vv��`��������o�WR�sѹ�x��@ykd��,22�&y��)�ᝨ�w~��T�6#�&�?=����>�P�}�!��~�<4&DVXg� I����]jy5���]� [���a�J]�'G�X""�;m̾�D/U��ߍi=����u��D��7�s�V�b֟HE`"�%���ȋb���0"�� ^b4�Nb�cI�0��a鍝�ۃ���N���	֍/�8�n+Q���	vf�{�o�8s�*����/��2��%)w�	���ǎ~',_#�Y�ԥ�2�C?0+��(�y�%�����qxhzSjikzY<���Z]09�pc�c�,��Ǽ�6̿:��sJADY��Ϩ���(���[ֺ�E����V1.���Dl���fb6꓁�fIE��y�	���lzT�h��!E*�x�7#�x_��t݆� W�U��+��̯�y�[ޤ�'l�3F���hc����ù��gf�ȣ�wC(���̔�s]c~P�&�;E�4�'�����C��xh�)f�d�	E�:�'��Iұ���9 ��XZ�%�;� 4�����h��v�?��}��C���GH�.����C��R1�T�L�vT�iwi�O���L�jMj���}�(|��S�u ��5?���
�d�M���#3��_vҎ^t��+�ծY�4Ӱq;?+�I˥�ʇ����ZV�>�E�0:�\�#%T0���?�CP�S:<��J&n�T������lM'$Y+���q4f�+0����m�����}�DQ77��S�iVdK'��kҔ2�e�\eS<~�~7e���q��9:(@.�<����*X���3�;+��0��sE���O����D ��L*#�iW�Ċ�Ja��$׼|�ޏ~�`#�og޶B�H�o��q�b7!�v�H��:SY?��Fc��v>��-ú|�ɗ4�I�0 ���*e��=L��fFD��"q(�~fя��vL��Ѝb�;XuQ\#�q��n�8U�p���;HӜ����dƢ�a �Q��aĄ���RGf/�w�
=�FK|֝|���)r�8:
��|����'fy Og̔oN<������1/�t�j5�<1R
�=UL�������s�=�jqŔ2ҽ��X�(~�N�_X!��>�.F�kֲ�㢆Nr�����B���\3M)H�@m�/�~�S:#:(���g�I4(�Үmi3�G���g�!������)_�R����ԡ��vH���b�VY�:�L\U��]��A�m]ʟ�5:]*�\Z8&�a����ySU�1��"Ԑ|ؼD�7Se�?/�����!��oD��P]�t���p�=�(w66͗ ���Vh�EP�ɀ��720����~��Z�5$��X��	�.^�!Y2���5���`AH�F�&��3���Rg��#�M�mH�ߑ�g��{?�6����EB���@���"�5��CL̻*Ȣs=Ø�E��y�j��z����5,6�7b�����Be)o�߀�lI/F�۶�dO�ܝ�{[bbU"�?���j�Gi�!_�#B&���l��B�_�:c���/��lR�6�E"���s��Cw1܃���Β��S�+g��G@Z���d��!OZ��ڑSF�t��}���_���G�0Ñ'5b]�Z��s~lr�4���Bm#5`��-����G}�������7@�:	
iU|IoYI��;��˷�W�ř��l1�W
��V�!�M�۾������?��0���j?d5��_^1ϻ�)!�C3�E�"T�x�JO[v�p%sH�����lM*��;�z��c�����j��P�d�)Wl4���=�+4@$�{���]��~˛��/u���2�.\�E���l�5ƮJ<��Ө�׫��j�4I�\��J����~���5C{���l�xMi˗LD�b8�Dl�AU����0 ����h ��S,9S��Ԏ��[������\J����$�=aWM%I��?WH��������e<�`���ȈD�~�2�J
�1h�*Z�k_���dQ�T���g������b���|3��x6b�=�:��D[�Lje8T��X�����'H����������7�; ��r��2�Z1t�7+�`��}�!ϳ�=�sJ��9�k����%��"!�	!9���r�O�/�΅]��r{��P�J.#.��z֜�4���n�v�-�O6
+d����}��$�ѵ������r�b9��1��#�J30�znY�E=��&,�� �	ڡ���:::��i���?�mɒ�.�&�fM��nr�a{����@�2����}����`ʹd�{�ni�����^�BC�:�6�ma�K��(��:��L�#	;.�,,��K�)1헰�z�JI�G��+����dc���c�4�k�7[�;KFm�����+i��?�!�37�wm��Nd����l��!8�>guE�oyO�y��֬aT]�P��r1���Z��βf��0���%��ڧ��R���=H�8	~��S��T��o���^�[��2���:7d�3��bCB9&���ڴ�ڰ���	/�5�b?mX�O���E�f�1��;y�Th�F+�~�ͱ=�Z��r�4��4U��������ؑ6C���9w�j���o��`5dٱ����PQ�C&s��K����$�E�d;wb�U�)���o��ij~�*�����C�'����k�[�e�fH������}�1��P��o떬(�$�����Z
����/m���'	�+��c�ጤ����6m^�?%��Cm���)�W�ҧ�-�:<^+ad�a%2zm1_�5�ӿ�W��b�4��xq
��|�4��n㏶�,D����`([�?��+��EA��xeۙE��^�sb�$�>]�z�W����O��S�y�ng@b�X�����2�
��$��؉�NO�������ne�=�&����wg�6�s.0t �2y�u��բZa�X��8Q�௾�ȶ2��5�TkAT*��g{��)� ~z��-7��م���y�w�^���a�2��D&fe�Mȹ�,�R��#���{�����1C�g�L�X��i�109��=���2�$4�Dc�
h�Y�[�w$&������m�l��)��W����%�y�u��_�a�R�����|S��%B+��u,�N6�:��x+��6�2@��U�þZ֔ք@��jI	����Z(�3�ߜb�*�Y�.�N�+gӘ�#dT�M��g{�{a�/N}�kʎ
MUN>��)�8J��Iv �J��D�s3qh!g���{�fX�c�Ƈ˒���P���$[����_��[�L%�O�Z�gsrd�p��5"��t$��\7�E� 쿓ג:��O�:u�밣�ػ�97����Z������T�d�3�ɢ+q3L ��Om�K�@����G�0K>�-B�*Cҵ^I��z?B"%�G�s"�r�;��7R	^J�n��3�ɞ����,�#4��/m��ۢ}
����.���ϒ|p�BNt�o�����ȯ,����C���J~.3�%q�v���1���5{��p�Bh��@w��I!!}h�om00wn���V��3����e*6=W� ���z�/���$	+%��yzGҖ10�P�^LX�D^0�y㝱��^�2�j4����!���ٹ&��)�kHf�XX&;���Ӻ���i�!٦`|m��D�+D���)Az��<�����fs�]�X��#��b (�ݍ ����9؈L�}h�M�� v���m������𢩏L̐^+\��?���p��}�ԛI���
���8�bk���$q1���R���}i��R�d�{r�w٥�K��ߜq�q%��¬�����9l`�7N�\�~�h���l/-}���{���Tv����0ts���*X����D���1��[���\aa��=O��ċ������aǐr��~w<��[��[���`��Z�(���Tj��㴚�������2E��[3���G�6Y4|�Eu;"4Cv��� G4�uC����EM�j�?}�����1H�g��E*���y
�6Xw>[ÕG(7�i�u�6����B�6�tH�Ⱥe�~��)�m,KU̿z�y8y���8�R.$�$�=3/��Fg�y�E�J����4@Y�����B��w;��`m���ɺ`�~�ob#%"�`�W��J#�p�N8O-a��V����`u��t����l�i��g�>X�����HO�Ѕ�L�ɡ�_<�燑��ka���*��D[`ԙYeY�˸p5�+XG b{�jҦ�	-��+��/&��ĵN�e���3,���%�K��-�г0�R�)�)SU+aQ����|m�X��m������O�yGY��_��.bfY����9%�(�+��3�yD0�YHh	`U +~����t"]_|,�oC�x˨�ץ���P�wk�Ѐh��c��Qb�f�B���F�]y���;NT�N�y8E)+ƺ����U���x]���#j��)�*D�,��]Cv2�V�O���6�5���"q�����rvZ�^)/�-+��bh=E K�m	*P��pr�<jܲ��B������3��K�Esa���t�ʣ�̼��7���`Ll%\h;�(�c'l9�X���d*���5b�� O�+�$"mW�d�m���UQ�'�U�$G�E��%��XK(S1�t�Y[I���Bn�
t٘�B����F(��=����0kB@èО��@C�uQ�L}�-��X �XD�SMS�ө+����5̅��g_;����I �<��#��IC��	�ߤ�"��eû��� ����K�[�8u���|w��ء��Ao�^
x���v�Ì�a|k�5Ք��7�1�B;�ʏ� ��t%.b[1��ȵ��!h�d��bSuk-�f�AG�HhL�Հ��W~���UT1�1�W��%�t� ���GY
�ލœ���r=Gٜ�[qm�.�R�� @���@a��.4�����֯\�ʷ
!a,Ò[����o֦ q4�<��k��S$G�^����,�� ��F$��` ��\�>F�E<v8c�}��>�g�r�Se���`NC�`d[{��b�6�Z�md-��T�����X�%߽%�&.Cн4&\aʯ��s����c�X77]�,�3�O,9��P;�j�6�ط���O�Ϻ�>�m����C�U���OЏ+��+!�2����O>����
_��w���ƦL=�/U�d�B
�X��U��o��JG&�nV;[��sğ�n���W4n�$r��&�_��c�hoc62�Q��n�fz�w����[s�ju��I�Bg8)�5��XzKDB:h�O��
�0pF�2KZ��:�Z�ɰ�bYyt��+���!��������%�;s4:��#s�q��y��Nj<`m@sH�i�0:Yl�?%�頰@?��LQ�`g���)kU_O%�E������>�r�E?���H� �S��ѧnq��}f���q� m�bJ�f�$^q�iVP�t��撔��!8pA:�Q��놇P�@�Nm @`����Z�DĮ�٪�R�2�����Ǝ����{.���:�(Z��a��a� G����S�#��mD�E���&��2mU�J��D����U��c]��u�0�t��/M��]�|��I��Ż�� �*Z=#�����Ӽ�w�D@hz�6������8�5�0tP�'m�i����p~&��2��FI(MJ������~DED�1R��h�Kj�cש�ĳ�u��&�M����E,ӹ��?V,`J҆Q~;?���C��E��(���;'䡩WT���wz',I�_]�omw?->�N�5��-���"��c��"�����7X�F�fq�,�/{�*���[�$�}Q��fm,DP4�M</�ު�$���`�:1���
���!�Z_���\�S��\;0��$K����^�R���d *`zQ��N��%�Oi�b@Ö�
b�Э�0�M���M������b#�s���Źi���v��,�^�!���vd���gv�绥W��>K�������yD�\�,������{ro�9����G/�m�b/�D�2jl&)��d�y��e;�~�6�?}��� M-�wz�W:�-��H
�. ���L?��+V.<^��g;~�A�����$�	��{�*���f��C#��Z���f��lF�_��r�e�-1y������ޖ���X1��ԗt ��;@��W ��ٛ�	<��X�$�B�`^ځ F��������h�5�	�Y��a����q�`�������L�χp�u��	5�� 
���L��X�f�^�үEy�����S�����ӆƙ���G"����|����O���BÕ@��r��B,?�ã�=J��E�KN�g��
�3��m���o�4��
8K�^�4<��P뷑@E�#3����3p�`g�x��o�d#k���=��6�FW�3�JTvM�'^����ç�(�&I2�g�|܆�CH�tC�LESJ�H�~X�D2%�q�E��
��7��nUE��G���w|'��� ���!��L� ����)z�_�I���Y!;(�٪�#۽9G��O�d�g;�d+d*�@��$�����^���]�ZY�g_�,H��Ŏ���Kى �b��eM��^J�q�[�P1��s��\/HDz���vs�3 Y�hT_�.o�5��S�q6�!�;��WT�-*.��u9�ɸ���e�L��gB�ɮR9�n��%�� F�L\:��R���Ɏ��-".��;����9
W/��"��E��-!x^��>��#���M����o�R}����
�r������Xk��<�Y��=��K�4�R����?��GQxVt�� ���r��{2zT|Y��;��`Q�)�u�e�Z}$[�&�$�7��"�/��K����{؃�̴�gX
���B`�Q}���Q��\[	C�_i�,%�1z�+}��%{����gr.fh��TLG	%+qc�[B�7�j�!Ѫ�>�5@D�a�ć��p�_ ؾ�̄�!�*l�Q���u���rk$�d��b��;hF./�(6���#_�$⻄����m��;�w���!־]��;��RX*���/j�դ%n}��b'2n"�:^�����:�rT)yq�)xN£d�'R�i����|�\OEWT�V<��5�vU
�A�'4�ӽ���z�nE��m[X4,���Ŵ�̄q�(1���]kj��ۺ-�Pq`(���Jм�)ޘ��WAۯ<�Sƛ1�`xe��/�'a��n�u�oO��q��r晗�����Q�U�z�����B7��'�nF�$!{'l���|힭�@9	�9]Yfo��١��Mh���bG��}�)����%7$X�~[�{%%�v����,���� &�*��E�E�NF��@�W�W�f)Q�K��	��4���>�m(�r��E Å7�_#�#f��U��IK�y�&àu�H�g��yԝ����9���m�L�!(>*�^V��E|�� ��ߞ(>�Jua釾����?{]/��h����d��|W�.ȇ��]p��2�t�S���u_��܏��g賦bi-W�@��<�:s__8fa��-��N7���+�P��L}N6n�NL���h���HӲ	�p��p��<L�<ɖu��*��'����d煚v�Ag9�]�P�M�b�d�)L P��fw�S���[���e���7��m�|q�e�f��̊�<t�����������yG���MB�neGB����CT_Kf0y���#�@#�N��>��`�kx³E>�=J��$U�QҰ���o�ZŇ�o)��t�k���q�*���7��B�T�E�̱��E��z�Ύ@� "�4fO9���h�p;f���e�4�@e�R�T#���}�6��»\��h��{IEni������T8�q�8th�5Lއq��ef�����[�&���{4�6�vZ���c1���Q�i>����6vm2�7#���~2�1���Q�zVPK��@&�[A8X󢏴i@���oH�YfmJ87��\/�gw�幡+�?Q���Q#���sjsm+�r(�Ǐ����-��7O�|l���ar.<�nΌ�]�����3,W���'�=f��u���~�<����֕nM Պ���m�H�8Bw��˘[�����|��;0�:~��D����VaO�Y{����1�#��1�#�,�����|���}7� Ev����)<ǩ
j���!�u/�.ߓ�sb�[ҒJ�t���%И�O.�,sgu2~&/En��Z�-����>8daŜ����:�@g�%{�ux�8����*&9�{E��dKɰ�_�Z@���^��_�x��6Oe'D����a�t�Cɏrē�����N�%�Z>���3�@~M��m�>���V)��-���⿔A��M��(������I�9�&׻f�y<����Q�QG['��X�6�"��?������#}��1�탱�W�L��ZF3��qtq1pD��R�k&����{���B�$g_�UE�#pA3�� ���1i��@$ �C�'m�	�����nʂ�;�̥*���0{"+������9~J$���7�������MC��LOÒ�<[��}����7��)�1�3sY�v�+7��n�0r�m�w!�[��c%�0F}�O �6(����8��R����1v�t�z�z�ꦵ+ʗ�6�Q.5��b�y/�I��7M�`1�_xed](؉����ݏC�"�g�q����a�L~�6�tHX�X�]�N��ЊD���(�s�z��3lqH�ͧ���c�U���_��>{��(��U�4T��D%.�cg|j|&��Qފ�4�����bNUM������CU�܋⏁~<��0�k�9PE_p;��1h4�iTN�c�������E �f��J#���>@6�n���,Φ=���Ha]���l�.z���;���-]��?�2���-Ȭ�ڞ8�!��a�D�X���ŗ"i�����)�{@-�"Z;#s9${��s�A(m����H�.+lE���.�X���ū߶�c��j��G�_�V�Ϫ}��E�p�5&���:./{'��uЯ�7ksAvF��O�b������Zt���(�4����y_��"�9D�ھ��t��ޓ�X,��ge�]�W��KH(6�ޡ�[�7ȑp�0�� q�2�vOI4����|���b� �E�V5�=]9�����K�'1������럶f�@O�A8c���D���\_��AzW.�>�L',Ϫ�F@�o�~b����p�"�Z�/t$-� ��8	��K:���Ӄ�87�Y϶Tt�P%'Aޱ������s^f�D.�pU	Zf�|�ƜFN�*"�Z���Gs6*�����G*>���t.?��xMmw�L�<��Ч&1�}P���٠w���:�������^n�E?��= �J�2�5�q���}չ=�c��k���据�T�Ri��X���8�����+��{�e�
���|��}��v��$���}J^�f���;��>b���w1�`R��K�Zm���TC������E����Ә�n��r�7��o�>��ʞHYm��)�H�����B q���*H���;���5��Q�6������v:o��^��<R�Tu,��h���E��w!�\7�P���y��r M����]ؐ~KG��Z�
U1,$���\xV,J����8���}?�*��_�V{T|G_����$l�1	�Ś/��P����CN!�*KG��¢[���'�4��k@�'�5�����So����/�MJ�!� (��k��`0�5੦��x�MO�ZV�' �.�%) ���I4=�>)Fh�xC�����C`ڴ3�w傅*);l���px� �k`n�Ii�X��IlQ���2��;���q�2�v�i9�rA ��``�Y��h��"#0���>q?B�u5I^W�#=�UT���:�\�!_=��H�����蜽�� #���a��ʘ��%�����>��:�j��_>�?�ᤊ5#��� O�P��0�v���;��o��{�Bҷ���^��A��4C�k���= ���S���5$��=�*7�B���fy6�gh���E�0c9�ķ4�Ȥ�7�O0/��@����rE�bL�`Є��w[l5�66�t�
�u�����?-�@�FƩ�p�wqk]�!�rtns��k�@W���x?�F��s�����x�nY��V=ݞHP��f=�4~vT0�_ʐ�������@I��*�rܕD�n���3$pvnP���Tr�ҁ�H��P;�G )O�LPx�-�-�x�j/�ۀX0�w��`�J'(�Xׂ0��q:��%���\�us�<�J���$<�j�nxzu�G��A�'����n.�LҝX|�K::��,Lk�f�-����^�B�I���:��25�ޛ�}�Rq�^��o��wx܉1@������T���琅 ���)�D@R�a�P�)0bǏc܌���Ȃ�޺�n峱�3/�_�p2
�*+s����25�-)7���aF�5�tF�{�;r�SNt'��<�K������Y����ݍu.��(���fյ1"����*}/5�����8�o�ǁ�~��~�y��@�2B��y3��	��Q
b0A�F���]���<ëFk�M3c�l����1G��9}����{�N��b{�~�̀hް������E���ќ�>|��[�b��7�o�3Lz��V��p@~���Z<QU����5U�^��<u��Դ�	C�`�(:�xҳβ�>�zI���]%�@mQk)�嚣TT7�7�os��,iQP�¨6�����M�4�s|eب��ä�����,�K���FM$w��o�3$"/Y!�`��aø�Ѳ�؃F�//��~�ā�� ��,3���G��!w�\�"�}�����S�yk2��3����BsCp?-�Y΀�������@�U�_���<l���fr"��'�r��X���>4�>�j��	��p�I(|�A�*S����ާr���~�m�XV~���oB���N���0���	8K�C��mLx�[�p��R��%bp!���z.J���{LV����������Md'
�������ȧ�8��+jc�ά�G;�D�L=���W�T'�~�uj]l�$��qO*��,�G6'���/�^�
O<��0t�@H�Eo�a�,q�穚�v�H�Ӈh'jK�>���"i���]K2K5��?/�����w�:TG�7��$�)݉���(���ܢ�q��/�dc�>������ ��a�N?�/�$��K�F~�������@�.ٯ�;3A�3�]+�3�����W}i�"�H�ڞ�y*dۀ����n+�,\tB|Y<�����M��>���oH�"t�<xM�B}*�Ә�*���K�/�dI9������K�"��P��0Nh�|&�7T�pa�(e9�69ຐEg����2�rR��c�C/���H�%=��׫��j�� mHT�.?��e�q��|���X���#��`_�⏃P.ϱ!-[�PV�"=�Á�͎Y��%y�����9T*�O����S��E"e���G�w�9cKꂡR?�� 0��!L�^��g��]z�eK����BV�r[x�.-�~,�K���z�'m?L+�-�p%��+|F�澝#�!X�{+�pzN&(��M�ޯN�/N��n@���j����|�1�Ԟ ��ۡp9L������F�[�%
�ɵ��!:�� w|�)�HR)�峿�ik.�O���~��'"��a�|{���^�N?�K�Q �b:�yA��o�+9v��
����v�3��3�H�C�m>�!ҪA��JЯU&�?�D���j<�F��ź��x�Y
Rۆ�!Zkb�8�=��__Z���#��7������<���uk�d�:����$�SI�p)�1�?i\1���7��'�����s^$
��aa���w�����>��h�#�y��7�o��nl�8J��C!�,��g�A�i��H]+��yq���eM��m\dZ��^C�~`�yW������a��C����ġE�����I�n��C|��C~6xA��*9ǻIl�{uGͮ�|ΰ|vx,;ی�]�� �b�d���N�L�Ԩ+3Ȳ�lJl)[nd�������_bi۲��o����g�S�ǶF/Bfi�Hu ��%�g4=c--�*1\)<w!��0&�͠AR�(�R<%Ħ#�D��: ퟙ��KB�H���v�������L��Mp`�5���T����d��BIN=����s�~Yr}�Pm7� }�ݷ���k�c�;���J�}�z��	G�a<u��{L�x�Q�c�����?�(~{�!�*�އ��m��M�VN�j�\v�/��ǣ���U'�$�wC�g�ң�<�ڠ�*��G����eu��1+���ȟ���-g�s�ޮ^����M+��l��D����#hf�x��kOߙ8Ty���� �S2�a�Zk���X�9 c��`ސ"�a�b�-#mzq����1�g���!���1+bR�����\�y�j�n��z6�+�?12 �t�恓7���E\e��(�5]dm�~�L0���}��#�8a��� x�w4"�I�d����x*��x�_�K�Ρ�tFw�chh9t��P��^+���qDrF�
ޭ�v��� ]� �1C�BܨA�%����M�yH���T���7/�����	�Ó�����Ӡ5�&Tqq��19���j|Z/'A-�2�֎�p��KβS�@��0,�����H}������=������'����.n�-t\ZVk�)��#%´E�G����b�ԏ�x=�ŴD|�0�mw%���m��8:�ZZ���U���M{o��7��D���_��܏sJ����LY�Wsg��1Rz}��M�9w����@{���ge��Yx:���$g	)Τ��HI�����N헏t�D��](�{���B��1}f��)����/��N�/�	����Y�]agA�<����nX�y�M^x�`@wcIɉˋ�X�tQ����|3�G���o$,�~�m2�A^��~���JX-_O�����{vpx��"7Sָ2�|�Ln�ڷb��P"�r8�tms\!lĐKp긠֏�w���D	l) �͜w>s.��X1��g��%�+&�.�t��¤�:�t6Z�����`�z$�t��=�쨺@e�.5�B��zQ]�[q:==��BʩfKS�ǒJUo����?H�%�e��C��{!U�u�?�y��C~��M����rw%�L�|�T��<m�Xj*��-��5vQ}&M� �*�n�}^�����8E�lI_��w�[�5�Y}�x��Y��Q��.�X��̔H�����]��Cu�}��s��dJ���\:o��F�{�N���[��8�ˎgH솃By�''a2}S�DD*O�11���Mj�>�ȁs����k�k�kY ��;FӷN�� �[�О�o�|/���`�	��^��v*�j��a��Т�Yj������M 94r5���SR4�uNW�z�B�j�n�)���\�M�Ь}u�B�����NXB\�DD�6����e5����s������2�	{�N��h�XF��	��.� EA�h�Ra�G��\�t�Y�����_l��w�~;U{#�e�'B���tǉ���U�|���M#Uӯs�(+*��8
q�C�J��V�Z]�^NO��vJ���V�:'!��#R�b�5ӢdH�D��ϻ�K͊��8�>즲9��T���
a�8��!�L�i����1�߬L(:���ͼ��Q��u����*����us��0n�o��`3~���b8ъhu�=��j-���;�=
�Ѽ�%���t��O0GT� �2|
4�J���`��:r���iJ]px��LкZ4"x)L��b��N���d��T�C�a9/9�bh��/��ٍQ���7{�a����,�}��U0`"�aF��{�A.�H��$2�B�>֜*K��p������&2�,�((<���C��զ>آ�)�N@��!oW�P��=U ?4&i���t��˓1Y[��G�\-n�����tt��-_J�~'����a�Ь�N�z=�H�AM����̉�p�mQ�^beoe=g��`d̈��k���^<̩�e)�.ک�Bk�3�4[G�|����:48g��S��Q�`"�Y�/����z�E�1�~��L_�ط�D��ܕ�i���5�!�1W���շ�}J�<u�_�zF�K #�
e�,Y��9�O?b� P��z�agW�Q�~�\�����:�J[c^���4�q�Χ��ol�{�7��	��ȯ�8tRj��7!.7��|Ps�LV1���K�X{N��$�{�t���K�l] �V*�Ϫ���|�8HK,�a����j+7B,����.{�kd�6�O$o�DLn�JM�]�;�篜t��]��/������6��VM&�'=EϘ{�,e�^�w��S���n��ܝն?i��s*�Iʊ]U�?Iۂ��D8��`���^�b�TK�r�b��x u�	��>�w&�|���վ�x�l��	ٯG��^�u|�#蘐��|r�X�՛QS���jUI���5�Rϒ�<&	�_4G�Ru2R�C6G!~yy�9�d�Vsi���!=���g4�J�ͱo
4�[
�M���9�����9�'E!<�ZB���k��f�'�N2����/+�58�:��I�>�ip�S�W,�i�y����PԳc��0U�8�Gn���y� eM`N}�ߖ���n)�~F��6��{�}2�	r�XR��8��P/����5����.ۈPzGf1�8�HZ2H��L�!�ؔ��BSݣ�#]��{*=�Z<`�]�+�v	:.�a��4��ʃ}`M��� �� ���)X��^Y���%��,�o�Θ�5J~�:��5�v�1��k�����p��f?[&r� VO7�j扩I�:���p\�+N�G4�X{"�/mc��Ql��qkL�:w(!�8�'1���+��<��l{�ۄi�`
���l�즘��8Hk�o�p�il%���R}�qs4u���ꍜ5��:�I�e�T����(h����-)�\���f�m5����o�K.亲��T=Yڇ(��TX[B5$�ƺ� qi�[$Y%:Ҽ�P0b�f
���{:&���)����,N���Վ�.-�4;���Ţ�7'݆�-�
P��M�zΝ>���7s�ɗZ���Z �P��T��3+]�]��yv��vq�Ʉ/�	��ه�Hk�`D`���z��ZX�yI�Q�X�\(p�Q�_b�ͮG��:�	(G���dq{�v�6�iP���Hc40#����p���p�0W���bCBL�DL��7��Lm9��+�WDX9���S�W����Kv�F��I_��G-}�-�~r��Z�x�j�y��'>Mu|���HzB�[�O�g��c�����\�ʙAFa�{�+-*�,9vc��D2zc/ܲ���y�Ϟi�MoゴN/�õ�_SǗ* �s�Ħq0�<�P/�o�WdӈoKa=��q�}��$�,wO*��\���kr�g�t����!��s��@�W�d�Hj)���D$lŃ��uW4�⏞�'�5��o [ې�z+'������k�����_Xi��/nB3���>b��ƍM��Eȡ=GOs�c�EԺ�9�Z���#@c^�ΌҞB8E��X����%�w*X]��	N�|� ���26��z�w��?����Z��@){H+��ژ�K�{����Ny���P�~���d��*���YaF�b�-���CVE�J�n=�.0�����oS�Z�fUá}q��s�R��Z������(�X��eK;Ǹ�Z�0L�,k��O�8��l[iΡj%ew��X��!�MRJ"խO+��C�&q|�Nnk����{d:��W�9bR�����p�OU���e(3���?��0Ź�JTz:���B` �˝`���%b9�mO'����͈$�K��r���v+��w2 �uv\!*��?}�۵��~WWS��a��s1#�1��ޢ<, ��j�-@��]o0u1���XO����u<�����S�l�O�~��1Y7�jiA�i���I���x�
�Y����)��¼n���kG�5bX�@�ݍ�w���}��2]����sƇ#�
eJ^ �89�.(hL����(���Ar+�ʓ��h���93|sڅ�)~d �96�&��!���y)|���kX�t�jėƦ��-Q�eHӚx�P�ӛ����g_®Ӣ�]DI*Ⴑ0C R�ę��W�)��T�/�������!x/�,�v@�d{�}���Nx��������Iu�c�o�ڙ��R��r�a�Q���_x��sb�/����9�=+�~�������E˽� �.Xm�ɢ/?0s�	�FC����U�&�ޞӇ�JP5.Ug��hG=_ݚ̙[O��F�����2��F,�[��'k�{�+��Q���'�N��
�5��G�3C^hJ��A��g��^�@���&�dZ���ܚ&/S�_���8ߴڂ�2N+6�����)ξ��G�G�ʞȥ���ˏW���ϵ��r�8A�x�S��v�L}�D9\)B$S��c�8��CI�7�p2�Ύ�
�3��9�_���<�b{Y�q�����ʻ��HtC��}��U_��<[�hYYv�#��!���0�!T_�h���;�����{�?�RUKn�D�Hr�0ƻ.'�H|��F����sK�����E�C-�����H���W���up^�帥��f9��-P����Y,Qi}��s��'��@C��t+s�P9o�Ȃ�Z>�a6�"��=G@A��d!�f����.���.�o�wy6����ryHc�p��#z��aB�%G�]�	�x��O�OE����M�_u�\�|�1��q��Dr���b����l��YҸ�(��J0�  A�c\�j��PB���M����N+-�aΉ�S7H[�U�+�_��6S��������.G��c���0�Dn� H��˴�I!���n�f��W]�Ʒ1.e�3��
"<���Ջ�Qⷻ�Y�U%	0t�Ә��Z3�[�J� V�#�����*=I[F�c�A�$/g�H��7ufuv�h���b��i�����x�&Q*^h�
��K<C���{�;���i�
E�"��ЏdW��i�Q`]�7�'�w�Q��W!7��/Z��R=f�P����9���WN�?������ּ��	����Ja؟����U
2���'A���˵�D8�PG�#�Xn��˯su�*��}�jǈ��=X)���`5���1	��lܡ R�렱�RAa��3�[��̶r�gd�?|]��e&MC�df϶l��I��BlBz�(�)�)M	�C87!�:|���Ϯ������B����`���:�����-������T+h!��9}0o��<i�H���*�'6Jpg\�OT��mgX��|
�Q&j�AGo���\l%�4��3/�cyx� �j��2b�,���xRc�B׺g��ѧ� �I���I��i���4�f'UgO��-o��u2Ӡf��;v�l�n�,s&�j������a��n�AS�^t�mn��O�V�uػ��F2�&7���P�,u1��H�V9h7=��.H Jm�K6��R�-gK�,Uf�m��̛6rC���-�/<�e���g� ���=�|A�@x�j;l�ͬ�~���ϔ6jf4B�����m���\ۮ^W�����&�I0�d���\3O�á��l��!�~�:���/���[$�a��uy�4��i1���!N�>�,��0k74���Z;���&�yɤ���_�R�f�(��V���0 �֠rOд�u�7��6)��&�7�VwG���G{�#�	(ZJ>_Ȗ�d�1Y��=z�]xa�KL[��	(����|�*���j����qE0l;ߗgv����t~r�_�;������k�_Qet ��SpA�Yl,$|O'� a�[,m����F�m��Y�
�9$jNBO��C���J+Y�b�%�k�o:�[@h��]�ĭ`���w���@�q~UɎ��^x����fK#�w�yx��QTd���o�]������2�	��^�����O(�� +���� �g�;��M~>���ҔH�ag�}���}a�ݵGqH"��m<���E�k���W`�:�.�[�=J�k��W9���ќH�P�[�dYN����Eja0����$t.p�΀�d';��)��U1�ш<g�X�J7�Α�Xr[�~��[t�8�nB7]@Lk��d�o�c�)�5��l1]a����+D׻���@�.��O���~W#C���u�P����8�SF��Q�~6�2L��M'�&���Pg�њq̓8S �>�$�5��9��f�U��E۱W�sY�'%��WX���2���7�˷����g���r�"��达	ALr���m���	t�eG�{�#	�2��E�K@�R�o�K�����+��)ۗ�٩����/�,G4�DiD\�V��n9���􋶺'�9�R.�5�5<�K�y�`�
PJ�|�IG��pn]��q���3�fMR�QW{�A��^yje��>.���u�rhjYi]t�e�X�y?Sh������١g̓�M�/VY�հ��xE8�*�4g��G��|���TɭL�I�Y\��Ⲥ�!��[}�.jG|O�~zu�G������LdᛇFұ���խC�Žb7O/��o�]$�cJ 1�� ��o�6�1}���o-�B[����+J���9��
�k}�0����B��;�N+��^K��,S�}�y��׳�|��z�Ĥ^��3�ǮJ�=5)o�'�.^ꪜg���g���4>�A�*��;�rIr����m��YPr�E��a;�w[Hٺ��bw�AA<���}� �G����$�l��� �9)���o�ka�KP�U�':<:M�;V�,���,l�Ct-�)���Ń9�c����5G��譺��?�ɼ	��(�{�OK���r���T��g� r$D]O���:��:�/JU��1�e������fV]����K�Yv��2��i��x�m(*0�zݒTe�l,�����[�sFݧ]��\lj��Z��f�y(.r�-5��b&Q �3���G��V�qPC�,rU>/յ@p�i)ֶ�h�)1��"�L}܋�PIp����K��|H�]��¿$x�3��¿��(��H+l���p���ezxH��s=�RW�/aP��{��D��!x���e�E��ő������*��ȷk���{���L6شp��y~����4���(� 	�V��D���=� ��z�/b��WX�z+�6�!��^�(�а�y�|���Cè�|P���]��7Ȥ�6���a�PN�J�@��$Ш�t�</�����
s($:,v�w��]ݎS���9�łj�7 _Vj��!���&]��L����h]��^���P�I>QO��W���qq��o:φ�^m[��Zpɒ���Q�P;���]�2-��A�!1��N�F��	��N��6��4�|p�"=خ5n���P�8S`\���Y����$��r���t�;�`CYQL��"7�j!��s'lL�P3�n=�� )�CH,��`Ԛ '�2����S��b�5��03?�.���L���.�<=���ckI��� '�&>�;�f���o�,��S��#}S�JI�@�[�MB>�P^��#$5mz��E��=eQ)Q�#��پuRB�|�G����^?h�G���n���VVt�a�=�OP~5�;#g�`X�r"�>��P�_uo�Lj%��)kI�A���y��ʨ"��'�s-���dfiD����I�ۥ�F>���>��򘓢:��=Xo���3L�3��~-�����JDG�m��k�?��R}�AoQ����C����~�*�:��*�[�4�즽�U� ��α���
��Q���eLWu	׉j�F�_1$��b^��%�0��ۙ���HZ�<�{{�\5�bz����M��
��m��a�ϲ�	W�97m�$��q�j������z�>�v\n��{L�Ə��o���4~�3_M+��Q3��Zs�˼$�)M���(�z����.xʠ B<{$ә���޺VAʈy'�m�W�Դo�ZU@A��(*�%f����O"{�I�*�i��>��H�9�k��{�p?I�[��|f�*�[Ĵ����X�Օr(�ǟ�sL�-F� �fw��Q/�����^�>yS�gp��JE{I��0cHV�=�4�Z#f%��+?��ݜ��犕6�c�+��w��@<����)��i�R��;�����a���c?��W��Ž/w�������E�1Bg��89���oO��h�Y�����C�� ,�7���AM{�(O�r-�u��3`��>4�v��!~3���1�d����Fv=�*[�J���8Zu������8�W�ߑ�J�Bn�khڔ��n�ָL-�)D�_���AX˯��-H��Y,��0[�_�v��qh��އ��N��Qzm=f칡���'?�"N��ɨE�����y�0�� Z��C}�W�-�F]��@J2%�(��J~d��5KNd/j
O��X�l#y��!e�v����M��.I_�FPr�ɮi���s�غgOZ:�J+�g�>ڠ�b=�20�P�����vLrK�G�S��ٞ6 Úuv-Y��i���s�&Ep/��G�4H�{��k�z���;B3�q��1�q�'��Q�7}�	{U�"܉�9Y�"η���o���h������@(����Q&���.>p�]�ܪ���D�q'�.5P.�ݏ��L��N���(����ф:Rҡ�̎q��C-�G3�B�@ͭ,�2�.�ő ���U�lE��̬�}����Ef�^Ia�Fw�.��wkkV��mJccp;e��]L�$����Hl?���Ul�,r�)A�)\�� 6Z�~�f�8�*����½��UX�ۚZ˱���>�y���s������I��  �ӾU�m*�M����aqdmf�b.Y���+(��5>�j�ѷN{��y!���&0 ����	Kf�熦Ŵ�(	��>��5�`~�,�<��p��O*�֓�_ce�yu�6�@*f�G����7��Sǃ�_�Қ0�$��,S; ��� ���Uc���a��"�_��v���gǺL|��b ��8��'1R�IFeǋ�A��	*�g9��&�����m�%��5j"cI���'R� ���z@�!��N�������fXߗ�.��n��:]:=�g�Ԥ�mBGYv����S� 1���X�P��f/�Dܿ3/��@�R�R�3B��g���;H��~2+Nևh���Ֆ��[�2k���A�W�����r �1m�:M]V(tInVV%K�z��c���_��IAS�v-E�v�����^�j�;��7�xz����cx�+m���B-�hF5w������%+L��/��ߴH>�l(�m�Ϳ�ԟ@�;Iq)�o�"�)�T����/U�R�߆�<��������6r/��J0pG����ާ4���a�^q�a( wFwk���*R�^��_�>�|���uG��i�j���{�s��]�̍ݪ�-��|��e�ف��秏��0���D@b���d�Y6e��?�2��ӻO���(�z�&d+ ����"���O1����4�<׼DwKB���ݷݝ�[b���j��Ȣ�?�VO�V�~�ZkXS�Z�=_:BSL}��G�	w��R��5^T��B�5iì1�,�S��}��q0��A����ZI���̲T���k�\�+Ӳ�4M�D���bx5~U�;����FF��8�]غ�g�ŀ�#�;Ѐm �*_���u��!��/x(�,@�t������}?
��@A������t
Rb���S�x����$��¿�.����p ��{�!=�qqN>ԛ�dOc|IKi3š��!���~+�UUH��(^A���`>b���#<������y|�Kl��KX���TԨ�A�8)<ƫE�E���(+t������������Eϔ���(,c�y!
�(*��_�Yj�?+a\-xJ�����!#�ߒa�~`�ܯ�
��j9�m�&׏5�E~��穘�yy���	k3���y�7� J�6F��i�ʙ~Nb)��M�%�� u�$$^ �e���ʹ1Y�yF�� |��I����W4;w���D�˵G��C`��:ik�P�� \�7m��zI�F}��oI�<�u\h*������ҿ�)�c������A ���RE����P%ɹ5*[M:8�4��+"ۭ @����5 ��6pATM.�&詉��)9�a�Qо��/|�1�0ͼ�Ԩ�h�0���3��0��0�,�Y	'���)
3�Ɔu�2�" �2P8Q�Xa3k^��κ�Q�$ȕZAE���sİ�0&�A�+��Bw_���̆��n����y�n��Ҟ ��-�s�5;��q�("iT��8�`���1�Cw��0e�LBuԠ6��ݚw���C�PA���fk�k�u��ۯ�`�sIEΔ>]4�3���� ��|���0ȕ3_��Ř4���L�E(4=�P�����x�}r,���	W��G1j��?,ʄ1gߖ+k�p����X�Ϣ��D��.Q�<��lJ\�RUtUX&fQ(6��r���|;j��)��S�{����X�����䰗m\P,yރ%�?z�8Y�i�K��j�B8ؘ��Tϙ_��E�)����+���-\��8�RQ�Q:�=�OJBń���#<'�з��&��%N�q��-��FW&�ǒ�������Z�I��U4D�	�A`a�C!:h#��Ķ���Ә<mE�<X��#����1j�{�NV&3���FQop�b{̍�!Q-^�:������|Y'OM�{&���R��~�U~��d��8�R��4��ǑtR+�n����C5i��ũ��yۆH ���O��}�b 0q�;�;�<W��'P�:�)���ě)ȰT|���N�jȾC*-�k�@�ҹ�K����I�}�M9��Vh�u�I��B�� f�y �'�gE�z�zk���4��/�u� �o�gW��{���G�F%��Zv� ��������ٰ���������k!�o]&U�fvI������H�7�����E��P7�|��ߣ���NX�f'׶�{�|����c�2a=�V0H�R�<{m��̑v
_p�X�9 ��!�ǈ���˃g�`��r�Є|���AM������$��Yѕ$Vu����tȠE0ѱci7�\�!�����o ���W����8�*���h����ʤ���C�:2#y���|�2e�zL>)�4@z���.�iV�۪?�%G��G�9EN�BH�ƝH7ڒ���o�����Q`�F
sY����aH���y����6�}h����%֨�k�,���N�)u�iNP�AC���ћ4EI�t������K����/
/.�kI�y���֐n��m���~��c��uK*���ڎ�ҏ��	<�"���_3�>��.�B�-�f������14� MMt�_`��N�v�dfv��c9��0]��Eܭ9M�E����_rp�.'w?*=���4�+ȥ]*�]�����ZS�%o�ǥy���q����I x��	��c�hҐ�FGnNX�V�N�H��`�Zp�r�@{������[3X;!�dkqZ���������(�<7[�~1����_�NZ3����z�����@|����R`D��X���}�Z;4�N����$M��}a"%�U2��:eȚ.����߯c�0�#q!ɛ�������؂�Ku�tT���A4ox����㪶a^d��'��MM���6��X���4f��y��W�FT.f��I�M� �R��z�TV,=E�K�� ���[p�F�~���_�_�)C�g},��x�Ikq>��4D�irL}ԓ,$����V=j�6�t�P�v��=N5�~��K&:X�¹��3��,��n*��e�߳�K�l���	g�c��&+���*#���K��i�������[;O~+0Ƕo�2���*C��5�d�N�!��0�,����l��Z�R���J�j�[�����n��~e�l��^�f�K<<�"�o��q<�z��J�y���QhxW~U������h�O�g�d>
iq�O��:���U��m�g�)9��	�x����c�h�r����q24�_):���DC��*��,c�������&������$D�/�H���M��VH��fҧ<X	�LE擣Hd��5�����ed2���cW]�l89_=1�~��_����2��4w��q���f��!r��){(���� w� �3Y�5�,ʔ:Xj	7e��vW{��Y$A�>��Lb�\�	�Vo���$<��̃�mNL
x����l����<�mu�哻��nM��m��=x����P�W���IB���=>� ;9롁SD-x���2,�F�Z�h[��ާ��-���4I�/C��,^�1�y�Fmoa0q�׀d\	��]~�M��~Ѫ&MB���������ұ���w�?Z͸k�Q�����J�!�1��2H����S�h��ryPs6`-��,�vd�C棞�:/H,_mWu�yɕ>/�~�_:�$�urEKw[��q�`و��ʲ,g�_��|j<|yb�ƠUhZ3��UMDI6]��� ����Pv\�1��8r0o�#��:@���h��lV�{�� � �!*`��&��I�k]�
�,ۻ����x�[\'c�J<Q� �'`{����|1Rx��z� �ѧ��U1�8!�:�Ld�R(ȩ3� �c����q1�8�,��nf%p��c�JY��#�h�1QD*m_h���Dd���<<�����ϭ���(�/_Vb�㚖����]�E�h;c�H�	h��1Z��\�~�Lf�c�v�Gh�u�81�|�?'�s߾;%����mN�yX������;�#pE�\8/!��pZ�c<�h�j�qG:%|"FD�4�vLg�l��C�ȼ̴Y�tO��A���uH�[�\uȨ�X�>I�AJ��ճ��Rx�e|���f����|_���o>�-x�s�?_����L��������6��?���5��0��:5H�	mV*/8b;�
�U�YOo^���5���cXԋ����z�Z�N6�nG3�����]�1;��3�Ѷ5�I�*�j��jP	v�	���T�d����
՘�ҟ�g1�NY������5������)�7PVF�Um�(�4}	39V	����%��?��Wuv�yCrY�&s��$��� �e�����Ǡ�����֒d�鶛ڛa)K6�J��i�x�_�_�`����������!w��5�e6���P����ofg��＃g63�Ǎ���↫��F=��',pB����B�3V�Do�O�&&3��I�HrJ���� �x�lܪ���s]��?����i���<�>�3�P
ۘ�}���[��P�jͷ�#�6��=3MV�Ԫkssϗ�>�u$�#�l����r�c��(�r�Qh�e�t�`��� �9� ��2C��=�e3#(��	�e	�"�%B`LG��Y-&����Ȁf���pV��n����w�I�� ��p�b�L��b#���:�2����&��XB���z�J��Niڛz^-dC�8ն��̊�K�rj���9� ������ӹ��{���fl$P���Fڷ[5#TaMX�{-=*A3�0%�kNӜ���h��='��������a5����(����y�x��I� Ҁ��=1��Q/#�9���v�fі].�6�I�hx��F�&~���Y�J�}U@�G>���uN=�XtQ=i]V-;)�GS\J���k�.�����Z�5H,d����";D���3G�x�04�B�����.�)���w�<G����:��.�H�nhd2�h¦)����}L�0.��N�NYׂ�X����ǘ!�����|��F�?ⷣ�a/w��o.<L��:�~
��Jl�E�0W��g�������>�Qr��9Q:���U�(�(��؇�ZG�Hz�Y00��?:�q"<��D]�):�90��=\��G
��#���|(�%={	���^l��v�N�G���**��"��`�r3�P��B ?���m�������Dh�~��L*�_����h���Yf�����E����V'��N�=��Gܼ�����b����4�Zͽa,�q����� TzjT7�HX��4�61���F���;��A<`�٪���,������2�n�N"w�����I7(�����L��9����R��:��P��V�њ�pR4�d^�����o�JŘ7�1ѣX�-,��tSe��ɮ��ș�2��=��Z���nHD�S8���Vw]"����}Ӝ</��&뱛�P�r>��qf�w�ݒ�N{M�&��詑g�f�^]�r����tE��	XMO9�t�N�a�}�
V_&�־��>Ӓ�].x���(
?&R�n=
}ǌ��)%Yݻ^l����=��p�	S��^�o
�]�e�R�TXF�|��^��ˁ��.���%),�	���-w�v�f����z�u+�����kO^W<>J"#��&�C�7��g&ԇ4I��0©~��|����^��&P�������0q$�/q"w�`m7�}��+4$FP��8���Q^���-�yCP���
<W9�x�^񚆴�$2Q/�^�U��M1�V���ӟ���X����2��ŎplE���e�΋3�/J�q�@ ��ٵ��[`=AC��KJ��3-���-�f��?Q��B��J|Ɂ�f�	e1̣�!J��~��
2����$�T�P�F���рk��r&NX�yDz��jw��ֈ���s�'� ���}�If̘O�I���z��CM�rT{J�J�&��᧘�nǈ����:��B��W a������x�}�[\0�� f;FC�ͮw9�d�e��%ĐC����9�����r�'�O*����w�,U� ��Ï�V�/\�G��\�n4IUu���B��yt��U�N�w��������0�{?(@h��$ü�t�\iC\9��I�.V�{�5�����z�+v�u�EeaI��]$���/M�Y��J0G7w�p�����z��@pDn����o������uO���~��Z༔'��wI|f��-�����H6���F��$��w!������Ws ���x�ar�i?��[�V,���"d�vDG�6b?�W�C4qIMej��oAnl���ɸ HC�&�Ӂ��r:]��J�p���)��S�DAL]@,\#�Ȓ��v��I��R��/襂F�ߴ
MO�E���Z�<�N�h��je�_oMlc��&����)~�n���w�G�1���H�1-��%'��"�s~d���~�QO�z������nނ?�y������p�O8���F�l(Ju�~�F�]���l�L�?ц /�O��<'}O1.�hKċU��Q"�p��B�H��ش�������z�9���T�+�cg�W�us�4����v�DYR@�����&9�gl=4
s(N�W2z
KB>x�d�K�hJ������\�1�f�b����~����;I�~���D3V�K�������-��dN�vv9O��]���񛣲�5�}�3��dE/����@��R�.����xV���jsE�!E\���.����a��ͷ%ݷ'�;2�� q��K�T�6��c8Y�P .�Z�5��;6/�Iylh��]s'Ж��>�3��D��1f[� 9<
e��!�!�7y�����O~���p���B
 <��W�'Mi5d7�Hdn�Ue:"�8ͮ��r���O�3�~�������{l6p5�4T��~9H���6RF�ζ�;S�F'�gK�B��X(�Ov�7���st��TF*,���$��{0
�A{�*ɕ��L� ��d� ��!�|Ә���ߌ*���V��\��
�y����E ��<���n��"H�7�`����_�9���𔐙����6!x9�H��|�,�ZCs�D��ahM�6n�]�4��/�RO�8lv��L�R ɒX�a�?Pȵ"Lc32/������������L0�Vf'']��s2-�c^�������:`Bl�HH�iB�>���1B�(Vzz��]@o����SlJ��:M��5�7���2��K�8y�r�]��mg�"�4��1��˰.�z�Ӡ���#�B�kx/�����)��5	,wD����=��Q�[Z�l�������f��ROU��cB=��֭���e���&e�֭#�ذ�w�������,Aw�����>�YR9I�{�n#�x�9*�R_��kH}[-��!4�k�{����rJcR�R��Q�4в5A��Gc����Yٔ^U^<�cG\`�x�%ؐ��X��/c����ti�f����"OIc����7_����Xfi�gA�ۂ )�*�[G�y�٬��-��ܤ��g��%m��8[���w/�6U)?^��Zk��*7��Q��o�x�
���g�M��ɫ���N�����P)�4�������Н�&��q�
\KaN�wO&�V�ݤ,+�IL�A��=�U��b�?.��a]�y2�.�
"|�1��f�^XF����9kGPt���)���gF�A*�ϥVj�-q�}f�L�άU�	E�f�b٦��,c��&:f[U���+��7Y��ԫ��9�����y�ƞC��M�d;^h�G�kS5�m{�l��y��Sy|5?���*UV�� H��K�eIs
}�(P��t]f�ώs'{���ͧ�
���v�����4�G;V�"�=��i�]`@S�_l*�^�/��e�O��9Y/�6�C�/���2�LA�1P�!��9�^�a5�w��
E�+��[�k �PBe¸<R��Ŀi^�u��#��*�K�j��UN���a�v�8�M����@1����#�rJw��X��.x�l��_
=#Uơ�ͭ��79����[�. ۋF���H��JV9c򳉘�#�zJ0H�)���X��R�n��?��r��7<����U,�_��A.�7������.wv>��/��+��ҹM����8�%,�}jЦ�!Mn��$]$)#|�G��"��'���B�_�)�8�hX�O�� Ǟ���Κ�I��M���Q*�*j܈��B�s�װU�bZӟkM�3�f���,ɂ�V)_�Ǎ��v�m:*k�v�U���r�P9�	&�T  ��*�ېo�&Md3ǎ.������9�k|��-^�F�N5�N��$�@�o�(��n��b����<f�2��i�	1���;_ǉ�|vʿ�lH��	�5�yl#�U��޸��[v�|!�_�b_F_Q)����>�����nL��=V�ͩk3�I��Y��3�w�}R�hG>��H���He�]i�-s���,ٽ�4�
T?�NT%��� n��/�j��И�����~��=s�
}0�I�g����M�1� ~��]��}��YN��ޗR�,ǵR�>Z�d�A��E z��Ĳ�ݥ!ٛ��n&G�#�rx��w �r��JDF�<:�hLk)���b���' �DL�bݯ�����t!��!0�nL��>��Kn��_�e�i�W;��&�̓��nr��S���4q�a[�K9#ǐ1�� �Hw�A�J���T�� ���5�*~e�T*,ɝ��S��QS����x���"�|^\�nΦ���*\�R�#k�Ly,�������ꅋ4!_�4'�Sa8�ޅv'�LÇ�=L;�~��0�,�՟Lg�%�Ib���G$Ɖ-w���އأn��m�	���	)"L)/q�%�~�"�6!�&�Kק����i��>�����I�{�u�c�H<�*[?�Y��D�;�1?,\�	s�"p�H�fp|� �$1NZͭd�+C�b����_r�j���+�Suc��g�ˠ��V�e�1{���mU�4R��WY�������Py��T���+�đ���� �/�۾B�]�m���H�ko�a#)�H-�G	�LJ�E�Z=��M�S�Э����8�~�XW�l�z���2��V#2ǟ�#UϮ�nn��X⍒�@�@�ΤS�{P^�Iт���*u��D��L����POQ*_S�H:�Տ�pM��d��'��鎽�i.�UO4L�yJ���#�WX�t�Pʘ���[�,8�w8��vԆ��y[�I�F�EQ�ƙ2^��&�>秓*W�}*���g��� ���j)Qտ�g�D�βO�x�O�ڦ�����N��V7\�t��{����Tڹ�LSd�u�d �`�w+{��aNS�:�$�^�����.`�p(�1���(�'�>����fu�WBr�bh�d�)]aa���_l7��H����w;��!x�x�=6Ǫ�[[�Ox��Bt��e�7�V�W�t�W,6j~�%��
X�Ma#o��V1Xj�|��&ncuk�ax8��,�y,�p�U=��8uYn�:?���ŀv?�"\���Aj��?��-�7l_��E�|��J��I���W꒗�Q��s�}#}O��I���[�3��J�q�V��ч��G�;4��S���N<7a�&��~.H,)�,���`��.?����H�@���?N�#߳���{ۚ��!����Z� !«�Rc�����s����؈9?7�*���y���D����j�-�B���@;2���^8
a�`�n�C.D�|�-�<h�;��AkH-1L>���l
D�>�5m�#�mp��<�v�_u^`�C,/C3�H�����N��% 8��+�r�6������;nQ˂����ļd8���v��A*FQ�(��i��� 8�5c I
@��m�e�4.x�}cLm��۶��es*�0��t����ﰰ�J}|~ʃ��t��#�Y�U����
48�3e�?�oS�<�k���q�跏v5�T����%�x��T�D�$$��)��6Ĺ�������5v#H��,H0	��mt���s��FD P��i�ƪ�*[��֑ g�41[sU���;z{�:�i��m&1AA����%���ͺ>����;+���$]T�h���5��1�50��jZ6eֲ_��F���|s�(�B+㮮k�� �0[�8H�i�����b"U��aC�Rb�(�%;�1s�u4*gli"GS�����n��5�
.%��H�g]'����!@k^��t�6�$D����6�Z�~�k��y���b�h�kN�������bD-6��ʰ�@6��;]а[3������:�h��/��r����a���O&v�!7���By�y����})1��S�˲��ј��oKX4��sn�,�e�¼�*�&��
�nC�GQ@�ԫ�v�앸�H��v�䗹�e�ɚF� Eͺ��^C�������8��	�8(&����x�,=��@4�~CM%�t���_�?�jىi
�Rظ��a�'��'}SW���z�j/���>�:��'K�o�\�RO�R��Z��~�
�hy�e?�N%V���2�B~Z�+���*�L����U(Ȥ˩�@����B�T� ��JV(����$Tze�����a�&�H����
�IPC������.y�׀9Q�<��b��q�.�R��V)��' 6U>�kG��q�x�,��6<���m�O�ǉ~��-7	��ݠ �$��v�]6Xkn2^��,�͔�g,ܥ�2bt�5�¶�W��ÍGIJp�Z^�k��o�2�鼼�[�5$��yx���~ߛP%(�B�V��O9�VҚ�K����~��p�&wI7w��H�T�fwy�����UFz�0�=x����z|�+vB�Ah9q�n �h��N��:�V���O�vP������x�{��U�!4��&���w&���,cM�'�'�	Ϛ�~�(Ò?�L|K�N�O,=?�.��(�����p��k���j����s]��u�7�`�waG ��x��M�i��չ�c��ٔݬ�s�^�|-��
l�[r��e�$��bh�Ebك����c�K\��R�E۽��������';�5�6�?��o%-�����+�y���	k�NpJ�C��S�w[k�ހ���%ρ�K��a*�p+r���X�œ��	��w���2��#�)D*�=�P[�@��|
�7��VMGb��/��\�����l���c�nz��B���XL�'5YQR�X�śg��P#��R��]yܨ8�6bH�Whѓ�sz��HF����Օ�_�|X�vL�Lc��F�(��y����J4GT^^�>��#��L�yP&x�&�R]T�
;���Sc�9e���^���`w��f;�`y�Ū�i�NH5�JY���+-cјȟ`���X�z�I��ꊶh�Þ�$!v;�$��7a3v2yD����z���.b�R�"����׬�݆��O�x �����BO]��1%x� Fʃ��B6w�&~�cJ+<ړy�e�*Aִ�<��^Q@e����̆G@���g��H�1��cc�P���8u��@YJw���ΞW�Wc�\�qRCɛ�2Y{z���̣u�ʟB�9�g�K����ox�-Ovل��]�fR3ꭟ�C=�T�pVcabEy�����z���6O��|�5�6����x/(�$юQ,ǰ�
5h�൙ k12Vy��>����\&�������Q�S�><G����E�H'ť���Y!Sv=�COx�<�/�F_O$��V�7W�n1��/,��}qBR�KUV02��j>�������h�N�Hd���-�������������w&�<�����߭ㅚn��ɩE{�'����Z��ăד��1ޑ����?�?R#^�u��)?�A��"�>������X�N��XsMn%�PqUO��%2T�crN��([����ʐ S��:�� J�bC�Ġ����z��^��:��5��!#̞�t��"I���/Yס���i����:������h��i�,��j�>��#�$jYB�dEXY��E7u�*-�_"N�=�˝~���� �g{-�,�.��$�(f
|�z��P�s��F>S�R�l�Tjn}z����˘��Q�}�:yNH_x.�{%Sv]�2����nc���q��ЪҤ��T����`<�a/dtVw��uX�kE��w��8���֡�؛�ex���[/���7��m�{<PZ�ҭpc{m�EG���6���2�����lQ�u��&2�h����C\mӖ�#����ObƠKآ>��7J���|�a.�����`��t)�Dw�&��3]<�I}��l��R���"�[c?��m�-�"�9��v���̰,���^��\Y�R(-⏕2��3E�?I5�� �e��\.���vz�3�4̱�w��wQT�,%A,=6FT�թ;"����L�n[%�� ��x3�I!�����(��g�Y̚�I&�mw��\�l=H���\t*�}o6>Wj��T�οm��H�<2f�7Qڬb�p0�
lw
R�H+����2���7�ΥCqH�#�����"��n���Az��F]s>�w���T��kJ��U���G��
���mά�{
ߍ�04�I�e���R0T�CF�xB�����m������
�ԬE�Ã+m�t�R:�Uz;��=B�Xns��G��sV#M
~'��&É>Z���r%5��i�.����C\lJě9}�Y%u�����5'f�F��0Z})f+��BD���O�j�j����!��8B��J7|*�ѣ�,f�fܘ� ����<^��8��_�^��s�`�`y�q{P�ц#A�-�4�b����ƾ$/�1r�_)+�`͍����D�SZ�oJ4űWo?����&�D��<:���=a��o�����X�u�:�����`Y��w��b���uw=]���E,7��>�H*�b��}�]�=�~v����P��\eT�@�~����2��U�@�)��Gm�H��ȸ���L�4���C����s4s����ǣ�v��} Ŋ�dc��͠L!��_'S��� �����p����R����tJl1��ępxfM�5�����%#q���X�!�$�AsnXY�?�oB�<z��4�)�lY�4��-^����ki���h����+j䬚�<}��=ۋ�$�����>��0e��c��_��p�;�x:W�	��mj��>v�4!�`���˹��p�]JJ��2!���g�H_�T�>��qk-~�дR}��8�w*U�g��û�x2�"<^�^���z�׻����A ���_����m�E��`c�[�ϊ����-­@Z�4T�ER���	����NR}y�q�B>�<��-tAQ���g�� zA�� ��q�2ggm}��z<ۥ�I��x���-!�"�:�B���I���8�Ҳ0��>�Ӻ2������b>�/8��MUN$S���
CԐ��U4���[��Յ�$�s?�7��]�zk�K�§�D}�C	]w"xa`�:lKAlp�_!p�����mW�X%o��&{&�/(�u`�n�^
������2��n��ŋ�f��\1��ޯókq���L�����ded��ՎW��ߕ�!� �:��V��\�x�q�+:
r�g>���=��w���~Z�Lt�����	�*ԬLC��j%H��(������/V[Q�B��Nڃm��S�z!���zN���Mh�T\�� ptvq�l�i���� x��Vޚ��İ6'e�SUE ���7:�pʋ~v �%Zd^���<��}Љ�S��m@MnF�۞��f��A�J�(�1U�����������[��M&���w�d��6ǵB!b^���=�;�*J��8�>Z)�h�R	���0Cz���E�m�B�*��R�v�ιB��K��6J^����^/��K�2r����=���p�\�����y��Č�I�����SL����GG�M�D��֥6:D��Y��2~[��D��8�47��ow[�U5	N�lh���F��|,�=�
���+��!��22��QYɘ#!US�h� ]/)�r�rd
�5��&z����W#����*�&�|�j�0�x�	_W��U��%p������a��,bZW�~����yDO�#�>�92''�����,#1	��t���C+b"q?������?��CO��,��=��ֺ����3A�w�(�j������e�aSS��Ǵ�2JEjw�`^���ax�����1|�w�K2q�	:ok3Ϣ�ⰻ�|����SҞ�峜ZL��;��k������p�3057ߓ�m�?w
q������&<"�� xDrE��ž�w*�W��)zJ�У0� ���ƚZu�b�
*��I!���uo�K��(b6��\��L�2���po�=���,�Ĉ����g�]�&LP���Q��.���o)�l�9㇞�ځ��:׋�A[�!�|� ��D���3��w����-�����Wd����Bӧ�οǬVm�Lo	�$H;����.�>�\^�f�k
q0�`&��â(ɽ�^�Oȹ�б������'z�evK��ޑ�7�!Yn���|=�r���m��Ow�Z�=�d
q�U��D������|��ξ���|�U+�����j��LN rʸF�<��
����žZ:��Hz
��2��C9��54Ѹ� �^6���P��,�Xq�V��Wcz6�Q�MVu�E�����3@38��x|��YU�m&|T��W��G|��AP�V{r�֌_*�3ho����I���7=��Xi6��-h`����3/�˦�ecW�j��QR��i�#]���#`���g!{f-e�!��� B��#|�Cx��wll��_D��]�d���7�t�U�q"���t�+'rO:e��N��u�4Mb�]d�޺���X�6Qd���sќ����t�e&t2MY�9�㉜ApՔ�%6��M�t+z�`���t(��k��|<͏��1��KD�����*4�$5 �b�T�>V2s�^����B>�*H6�#+��Og�Dh]���)�@���{N����IL��gI��
��-w�(�R��	���)�m����A��8^����U��#Ff)K��N���*��K}K|�]��M7_��(]Z��O��� ��D�*s!��$��2�Lv�G�݌���~O��Af��x9�[��2�	���w�-b��:�s��~0pB/JD���\V�h<Ѭ@h.�lX~�s�&V��A:f��T��fv�8�%�xd��%��4Mˍ̃��r��H�`6i��IJ���CB���1� }��̶S�/�eU�a>����]�h�ʓ�z�=S�8&@YRl�3�ց/�3��,�m��M2��$��w��ά�/�dM�݅>�(d� Ի��$=C�fPL|��jr?�Fv7Di�����	��Rb�-
S!�����(�z��&��x�-�H8[��z����q���Y��Gł?�<����I��f_l�T��!���-�o��k�i����Y��gF�R�"��ZI��n��^�lI{��d�J^
LNa.w)&�m�ea�>33�Le$���?DV����e~M��1Qі4D�r>**5�k��[�o�$܆�4���pvU��ȹf��>���;uar���Ȉ�|aO8��qHB��<D^cߛ��Guꑧ���0n$MD��@e��/�=IXwtIa2Z�{�ޜ��:B�T��8z���f�T=��ۍX�e��eO�����B�ʃ�#��Ƈ�����ns=ECۘGɊŶfk�̋j�w�����ݗ���i�hd��bȴ��E˰�e�?��N�AѼ-�<���o��o���tCD_�ckI��F�si��;Tgլ
�کsI$�C^��;�Iz�v%�6*��K�]X	�!ĕՍ<4����R���40�33��DHȚx%���+�lz\_GH]럷H��5@[Du��b9Z�ٔ�*`sĒ���Y냸����){s�><��҈R E���|�[E�m bw��.'�rղ:�^�)�E�"��X<���}3b�+�X0$?��G�e;�(��d�<�ڑW�qT����X��vpn�MN�|���ɹ�=i_�A8�5gk�!:���"��C�������V p	IE�V�^Z�[�|��{��x�|V쵹���'!��[�pv�[�u��1 g8�J��{dm}��<���T"!�Pg�����
��mH�-�����h<}?�<�db"�	�6@���6ހ.�hmz�QF��@4o��mX�0�Sbx�#���TЌY1�	�t��UmO��[}�dT䋚��e��J�η8�2m��;b��S8=#_��8[6M��O��WGY��u�)}���w�՝�I�`JW-�{B]9(W�o�7�Kz��.�UT�@(x�	�	k�EL�6m;�<.��[d��b���5SD�B�A6q�����b��sQ0�?1�����vح����@|�_��.���D�"9~�.H��8�t]�^�`�[+�P~yX�Ix�6��09�܍��P<���5{�>m����K�V�j��V��A���0Ns�J��� ��3�O�S h@�����X3N#���KZ¾����'< �s��m:��7�K�%a��"�cl�\��;��Y7�%ؤU�i�c��[c�\�����e��0�v<����>C[��J�z�+Q�1��'�5�D�z�����8�C<m������zx��'��`w��1�h6p����O��ϔ	��Z�X	�?������~ڵ�d7��ŒR�S�w�n����ՠ��A�4�>Xt�[9����ʲ���N��c����s�Ώc�yۢmR�"ٝ>/x�א�J�˖����
iR�j`�lȅl��l��
N�i�i�-]��a��D�L�����|Iަ)Et/�M�c���6������E�$s눀��fH��'�BL?�`��)R�*��rA�C�TR|�n�Bn:�=!R�H&b�>���gmW��/��`�L��P�-�Δꂋ�/���/�0e�u�rk�.���H�ܾ%�N�B����'�UKۖ \q���LQ����6��������G�6����vz>p1m.D|�zME[�!1�  j��'�[\�����͖*Ϭ&�_���^�?���g���[�� mw�d�'v*�#&y�:S)���(��/�ٌTua�~�ޡ�գ�Zu����юycN{�E���5�V�G"��U,.�8�4u�����W\%q��}-t�4/�Oubf��My��L#��j<d�� Ii>ɦ�sU� ��U]�}����Z_�����ES������5�([m��d��8��p��˫����'�����}��`X��KzD[S�B�SCщ߿�u�f3`��;��F�b����(���lA����1��5���h�^�y�:�mFΦ�˲�i��̥�d{f��2�O��ξ���ږ/43Br.�V�, N��.cD�J�"�3�f��T3��ˡ|l�lK�N��I����Fu�hf���'+,o���_�@ZQ�0�s(��^o]x=�=�Hw�bO�c�u�T��۝Xۡ����874{L��~0�9	���_Z��ٶ�G�M]��s��Oȡ��W�	�,)%�L$��<�I�����<t׈0h%��%�sX���ؕ��gTb�-P�͞j(C�ҁ�������J<��榇��տ�4x�ּ�A��ӏ��P�)uL��O�pd�;H��^W.$��Հ}��=O�%J���9<W���E�7���/����n>�.熫s� �űű�t�~%��<1>�������O��%]�����$��R&�*��;ۊ�\O���G)f�"�o:嶘	�v��6�qsUo�.�5`<=�:�EN�� �D{����i,ݭ]r^�ٌ�cPS~��"��g�8&ϲ�Bg˷eնǬ�	����i���ߜ��J�x�c;�y9{���Wҙ����IVU���h�-����^}��Y#����[e}.�����U;��<݆�#�uO@���g�h|Pc�K�[.2mL����LT����]�ͬ��(�wD�y3�ȡ1����+��ݜ���`[���ݱ|F�O��k�o��@1R;���7�p���s(�E&��@��=adGX'A
���-�Zx��	�uEJ��i8���Z�+��ݡ�p-�f���^*	~oO��,�jT��%����aj� ��
��]R��JMy��>$v�m��<_��Δ��{����p�T+v|�ApB���r��s��Z%�I��6"o�>v�1.;u�bm������] Ҥ<O�� ���|>��IƖ\�@m&�n��To��V@��|q���x ��'&��JLOt�o1ѯ7�N`� U�(C;�=�5Ks���_���RFhY>��b�G!��]�{�! "���~y�M��YM�֊��WZ���\�5Ɍ㐁����R��/�6��{��Kܛ)�3����I|��gE��g���|���H���e�����X�Y�bw��e���ߑ��ĒT]��Ci�6{�pܡ����m٘�a�����nҁS���XÌw�yogc���qҘ�cIW�(�F�d�+�9��#�/ qC�+��E�?���le�#]:;H�o�%��0�_�Ͳn�u\�)vj�yVJ�0��L�Ⱦ?7F�8����H�0��5wZʔ$[k ��e�x�_��$!Ծ@��i�gt75����J�lSN�`ۑ!�vXPW�XAJ!j���
?�>�PK����Z�J���'�!����aԂ���p&�7�����@:c�2��L�^	\�-��;[��i��'6LI�?�Z��E�f[x�zL����?�i=�as��t̤A��$��AYzP Z�g ���7��Q��i�����v��I���ڷ|-K����"���/k�"������Q���E�����P�H_�2<�?�4��U�k�f#�%3�B�[���Z*��k�|EY��K�S\G�z�~��ƾ�ڧBA��_���*���]�<)��z� ��O�Z�1�{k�e�}�}��"�y�1Ԗ�����R��yzt�[� A�5�݉t���d+&ZU��Hᐞ_��5���w�`������e��u0��#aS �E,������sm����bޤ?���N@�OX�uҍU��5� �ak!Ho%�^7�_�!��QӃ�n�����!��6�<���DE����1�v�P"�K�3�����X��$��:*ǳ����n=5���PM=Q��}Ю�`ANDv�� �Y VGJ;��OX~F��ݢ�ˁ��_��f�ڐ�ɹ}�̆����L��ld�j�(�b̿v��Ң��xv��GH���+؄F��H�(n���ժw7��X &boO�m㭎�	OD����:D�0�-�"{+�X�i2u|8�W���*��|�v����c{��	tXǰ�rB00)KQt��&����w�����fh�@
1*Y�GJ�(UQ	6�>d�@c+��B��
d��z�\��}9ȝEw�!����9~�3����[�]#�R�X�#+u�{z0
�Kש��#�Q�`c��eދ*� �T�d�Hb��w�K�����x����)����C*�s�c$��iwb|-1�'!�~eY�Fe(�x� ܫP�4jn����/�g��[���da�M9�K����;����=����&�.����pB��4��Z4�<Soo�}E@Ǩt|.><����ڥ����ۼ�-��B
�=Ux~���2=VA.έ�j�7�S_	K�O�@�a�l���MvW�Sƨ�`z!��	�� o���3<������ǃӦO��AF,X'& ����.���+O��>�mB��b4b���xyR���s��ꀃu�.Hh�Ժ��d��EK8��	�"��xP2^�MvC� 	t�~�����)�ƃ~z{o?��n��V�Q\ 7]����W��t����x,�.8 �k��Z8�g�*�9'����

�Y
�HcA�o��%�e�J�/^��o/�6?M���I%O���u�q��*R)��&�/Q	�
��(��%������P�&q��d�N�YhPN][D=dB�x�M��`�ݨ���q���"��^iz�46d�2�,��Z��Hb��i2G�/��\C�y�;����B,4���s��v��*���̨��
i'�t�c�U���c�Jw=*hE��m�6=�_��J�ܖ,���b�b@�4
�]� �h?�]���7� |k �����v~pc�5��-���x�6ґh2�s-&o�ڈ^^���{DJ$�^N��@�+�b�Ƽ% ���	�#në,^�y஍3U�%�tס	.�(��0���F:�
ʠ�ܿbk��b�+� ��OD,)}�(f�;h$�Yr,~�U�W\��:��(�
��g�<BI�a銽�~_ <L>�<��"Lu~{�Gv��C ��=���.�mA��i���H�����߼n�����b=.	�����NPu2��r�bՈ���h{!>�_�*f��"xj\X� �{)� 
�6 ��V�~h_��U�c�mR����$�s�����fE/ &�;H�C���)8��␃ݒ�Qa\;h&SeW��_Q�B6L�0��Q�%f�3����d]!}�"M��!/U���մ;�\&:YU%���!CaN��6~�]jl��,�����%hR7Q�_Rt�sle�1�k��6>\�G�w42�̫��f\TYp2i�ۍů��5������`D�y������Z�D�=�]W��(7����)���hW��<z���u��J�����iza�{�v���&aiL�@uy�0k�]���(G	~�9
9���u��Zj����1eQG��nny|o7
Ï�h���}����!�`i�7Z�"S3��R��>&Uʔ^��w�7�<������;��}��8�t3Av�1|%��|���/ܟ�m��O�X�����;��!_���#+��؀a���L�#X���h�c(�����hȪ�����!	k�Z���^�j�o����Ah�k����x���|��p�a��K?��_4E�	d�� ID����#�m� ��;Wf�'�����t��d���w��K��x<��UƱ���z���������+�����;r<�%����'EPI�N�n�b���c+�ob#d��
����:�H��E֙ze��R�j_�=�p$��&I��ʹ���G|�Ls<��yq��Ayn��K���:��u2����8�ir����]t~%2([<a��톯�$.����E���@�V'������39�摬;nL	�lK��#��	�G�2S�;h��Y��v���.̞oEt��/�I)�+g�XBIU�w5z��,�¬z
���;��z�9+Ae4
N �G�����d(�A�&f,MZ��zVe�X�	{���ŐEGBe;9�0�`g=�^�E�5����(  �#�����ʃ�6�'?�=��ʺ��uA�ƲR�a˗-����{Zd��!{PFk��񆎱"a阚� Jf7�ً��b���W�ٱQ0s �6����g�8�u�2_�,S��.�Oq�\	���<�4���*Ǵ�g�ؽ��W����pTr�Rit�΄��H�|��������4�͂p����B"*�C.'\$��z��#�e��'؛ڱd����{�������!Qx�;O��,�!` #�l�a�`m�<O�s��~&����3�0L8�Lw�]p�����Z��Vz���>���� yz��E?��"g��/����"w�lH�K��_\=L�CG�{��"�K��&P�Hї\�ڊ7Z;zPM}����x1����x��@9�U�H1�Ǣ��K�HT������.��&tu���=��AHi/kә�Z]��}��Ɍ�R�����.�s�{�Hp�+r<W����BA������r-�/��X.�����T�vU�g�Vpz�͗/I���c��X#a���N�cx3lV�7l��5?��`��g�G�J�=�-*�)��q�GCLx6>�2�fD�B� ا@Ubwi���Y����Z��rE@*��Z(��d�y&I�2�7��=Ԕm;����Y�8��v����x;�3?���t��*PI�4C�����G�&},�>�Zq�`<�}��������J<�Mx����x'W6���z�^Pǔ�9a���/�t�;���~�&K�*]���:K;Y%����VP?�^M�O �ί�#�\h��*���>�8?|�|�0�����`�N+�ٯ���}ө��P�|�O륏�tk��(��+6��U�v�>{���Nf��^�󉿴�-�䅱殈 U���n��2�gi��S� ���O�|n�j�졕h�������J!�O�P�w6���w��1�w�I��R@���0��1D�ӵav3���a���*���`�Y��9^`BÉڸ�8�иP����&��`��ʨ�7�Ū�niR�P�N�tWg�]�[d���CnN|��sfp�������ԼY�M��p�(�R]8��φ2Ϛ|�c�X�X���Q)������� �V�)Gs����)HN&Q,�|�ىx(&YK>��o�nZ���b.��'ǯ�|I�GӅ�/��E/��2ufg_��wk��?��:Q�Y['W
M������[_�`�V�TmbP���!��i������*����n��	���O(6*��]s.4�Y	��o��DP��?�>�EY�q�$⩰��.���`�K�Q�����!-�5����i����ŭʽi���%[�c���C������_x<1�f�Vdݨb12Щ���r���������.�|ʌ_㓭�ʑߍ����b=��7��P
�~W�H来8ȋ�}����&�ՠ��͓ V���[S�S����X��)?M���Ag���y����/�J�<�nB�M�X��!�kJMZP�1��?j_���#��rQI�u�w�1eZ�3�|�2Lq�Y�vs��-�ֶ�V����HSkLC���Z�W�6�w�0^�dF�J�]Fd�,��Ǹ$�WF��_ޝ\���Fw�U\�aH��O%��J `2��KP���\㊢���>(�V�O[�,�5Π�e���;;�sx������l=Ӆ&נa>�͓x��#�"8-C��JC����?��NW%�N��9�r}��5*��`/���ѭ�ڶ���G����O�P�<��`Փ�x�-��v�6��Z�Mosw�n{*Ϊ(��f`k�,2�0Zb�X���^�K�t.�}�И���E�Mڤ�c���|,�@���h�����L��Q�����H���^��K���0>g��2��g����P�<$]?��%M�o7�sX��@��ލ���:JY�v�Y�e*�YS�ZZ�3�r/��L믳����{)A:��Sn�C"�ZD�x�F�ҿ�vJ�Ḵ��� g!yo�D� A�ۂ۫�@�&�6|�%�yZ)��[�"V�$$�'%�إ��IN���YC�'O�\}���U�:3m����k.Pn���m��]@wy��>�����2ٿRsK�%	AXZVť�ѢL��̓P@|��8v9���Dr������߹�ϰt ����׬���iG�фs;.'*�p��L(sh��]�8p�]������ǜu����C���L
�0������+`�:�h��{U6 ��>e������r�;O��{�<�x���:o>��\Ö�ď,���6>�>f�o�}yi�o�.[e�׻n���C� ̕mg��	�)��k�/��Q���U��C�<G�IlDߎ��N�㡑Z��9�T�L��F,$q��F�|�4�Î���<��j~�Bv�B��I��]�cZ�4�y��+�B�:��O֡��?��Bk�.�0�E�7ײ�9J�D�8t|���S��-��aq��d�wM�h�?��L�F���!�1Ѳ�S2E�����O�I����^�3�E؍�4wa�����oU]FS�rugkʀmںb���|���I�4�U����L��ܛ8�z�x�eVg����2��>y-�W��}з(��O�_���*�V6�����W燰� �6Μ��_��h�&i�.��L��e�46�'��L����ýR�n,x�[�&a�4�lɷ/���$���b�*���Ir5B��Dr���}G�߁.����rF*ww�7�L�'F ���`N��'2�[�s2ڽ _1�"K���0�!�BmI���WZ8�/u��L'�œT`j���Y鈭�F�E��+�;T����u���q|�#~>)���p�m���&�����\��ݾ�0�%�������ڕ��~U�+ٶP�\%�;h�z�Y<E��63��,��=�GAr�y�)U��+��t�Q��8�ދհ���"����b�ɼ�=�?�W��ܗL�R}�N6�⟫������^{��(��Ц@�s�^ߟ�I.��%��@�}Y�@�+�h���q���$����G�9�YoI��1�Ҍ��'�-y��I;�axpR��e[٢�OF	uO��D�n�}	-�}�P�`<�xgi\��Z;���m��@t�~p��
�Kے�JF]�<?F�4�|����w<R��|șR����)'�C�}r�q�a��_	\mS�b��E�@�H)4�Ho,�n�;y�.2�t~Y�q�ϲk� �R�0���M�������D
گ�h�@;�9%{��\s?F�asU����/�iW��QW�-��y0፞�uID�Fy�x>�@�B�ĸ�om�6>'R��}/
fM���q�]S����Q򛊶�lOY�Ѩ��T/>�"Wm���_��L�����`ڣ��E`����ϙ�.k~ "�����W�2m���n%�<���ֺp"3[G�Dܔ��f/��웱7���N����w��h���F�~NFx�1�b��7��J�ծ��=D�Hʧ�6�F儫A��0�p�'�cQ�O���Ms�s�߳����yud�j':�,���m��Ӎ��("J%�/[�UJ�:c?�S�]��s�6s�܁����QNH�|0�hD@�����o�y��Zb�gg����Iq5�7����*�Sv����Uv��ǌJ!�� �����F0���Z4���A��\��؇Į�A�[�AL����|	��J�z)":���D��,�r"��� ������%��K���������% S6�\��'���wXMԟ4FâKϑ�D�1��X�e�{��[��3�����uLP5L�b�_(v�|%�ߛ��������28��������pؓF����w�[��\�Ӏ����t��o E蔘��6��ߜ]1T�z�l����ں#K��n'�vx�,��ޠ"y���������R|K4��\�Лh]�xy�ǎ����� �Y�d���̚�o�BsQ���56�6�)��B)%Q��i+�D��ꗬ�%UХʧ�C��Η����h{��ؑ���Ar���5 T�_5%�<Nd�.�.^����48:��Ƌ�j���D;��y�*fh���!⼃x7R����;����dAp9�U6U��å�/O�<i��i��sb��B�^�'����l���	"P�`��9�?����W@1��%z��P�63"�	6c��S,Q�SM3n�e��V����@qw��*�02A-���t3�ؤkd򼛋�@2hE����W+�KR�eG4m�A��E����W�_�Iȵ�)���_�nn���x�&�>���Y@��2�'Y�z�A�^0)�W�Zr(z-���?6�M�o��X�j��%��S��F*W��U�?����J���Z��^�R&���~e��s�.�N$ z!5���H�C���jp
���% N��/�y:�p/ħ}�r��G9WC��`Ҷ>�:�i�(خ��o��Z��'����ޓ��#��{��Y@� Ag)��=�<�[��ȯVs']4��I���
��BK(���h)L�F@�>��I)K �wەS�4]�j���=��5WiY�ˆ�1!�*��"��"�su,������F��a_*O+ύw.Q��Eֿ��.�]��2j,�\^D;O�Ǳi0r�¿s�%؛o��H��Ĝߢ@����Q�&�ã}�f Z�����y��s���4
N��1�DDy혤�:6�`#�Q��י�G(g|�b�ng��$BD�����q㠎pT�w=t3�1��5X�+y���g�溔5u�Ԛ*>�N���De����|���!���d8C{�,˺�Ƒ]��2?vZ�� ���#���Q�|�.K���)P���݌v���kh�c��5��͘E�
���H�҈g�~BL�Ĉ���9�~+��[gN����\�V,��t���:@)�Q�R��/�Nux��c�.�L�+�[?iD��t$����8����@0~y������n��"q�b}�!��[ao�c?PX�/&����`�>�k�����V2C"��������Kh��!nrU�L46���v-�}τ�J��h����E=�������<��ʣ`-�@�E�PCt.}<D�P6+�;--���"�0su��M}������g��+O���nҎ�HYՀ����O.�+�������3.L� ��i� ���34������~���Tb5iq-�$�ϫ��A4�f�H��0j�_����Ԕb�0�zWwxuH�Z�]�sm�f�(�kw��7�յ;���S�et�ZJ
l���Q�U!����5Ӱy��UΨL��'�i���1(�OZ*ʙ����@�#�}Hu0�h�`�Ne�HƘ���Rk`�%��U =}��팍\+y��~���6��
�+�P%Ŝ���<�ѣό"�7w.a2����F����y�+�IX)C{��,),��B6��.�_���vb*Xk\�P��GD!\ �M�x~̋dկ�'�	'h�-�,��V`m��ҨP!%����ê���Y��U����� �:��\��h������+���%>|�&	�-����]�FT���=)���~z^�q�U�t�^p���{L_e꟯�Hz�o; ` Ȝŧse};%�pv���U���@[)�'>�G10B����bڛ�����3tJ�T2N����oݷd��1W���Q@L��S:��-�X�)��g�z�<A�� ���.��B\r�E6q���&?���H�82�c=Gė�n��J�����fA�3��#�J4/,u
��?\�巗!"��5�0����U�
�́�C0�Y�YTuK���+h_ի���T�5�8�������Y�V�ކ}ןx4<U����w�P��<�K�l��e9����d�Ä�I�y4K��D�҂<��� ;EC�P�y��"�氐{%4o��ޕ�<��1J.�7��Q~Bk 5\���1]HhA�b������ѦS�%��bs���C��9Q�:�-l�4�t����:��i���]c�[��&L��z*c��ʝ�)��� ��������?%|cp�*�j%2`�����d�����e�@��y�q�j�񎊵���؇�-Gz��.����eK�jۄG�c D�i�N�v#����*KzB��VF�S�:N�A���~]޼�ZjvgQ粻�����?��b��#�ͱ���=0ľ� x{�����+,g_!�k������i��ee��.��ɯ��bt�a�	�dj��΃P����Ƴ�o�NO��a���H���47�4"+�Ñ���A`q�ؾ��/ic�o��=m�)TƤ/r����P�^\��N�^��o.���-�K�Ң#0��r9�I�B�h��F)�.7��׆��f�P6����8�O�X2�R��(��Bye�Z@�[��P�ݢ�/��.��HŻN���\�V���4��g�@��o����l�8�R3bB���/:$ث���8�C?&�q�~�?"��(�p��/zx���$�4��|R�
?�co`dH����P��O��dʷ]����W!�Gk����(z.'Y�����ܓ�~��9Wi�D�zD��'�'�6��>��a p�����p��AH=?�Y)^�z2���S6U,縲�x����=ד>F�S�9#��KpM�����T~
n|�.��oH�o���ӿ�Z{�>�A���շ�|�� $�CN��+�ض�}�����]�
�0��tn٢Ѐ�=��n��i{��3�aFwY�Zk��dI�^����noƷĚ��`����������wFʛ+Y�sHk����i�~[g�Ֆ��ŞA�$��!y�(-�^[M��U�d���N�w$6���Q���A�x��4��x�/8Q�S��=>��$��!dm�!R�S<��<�U^+0sWp� HV�Q-��2�!~�K	$����8����BEʋ���8�^����K��sӶ�����:���ꤞ�5xT1t�^T��ݛ:���XTU%�������T8ѪRbv����{����֌>�|-`Z��y��3�z�6Bl@]�y�@�?=�g�3Q5L�﮺�[+X �a	p���������R�n�NP��"n�@����}�f~��x������{��0@�b�U|���X(�'ٽG�b6[��y78�s�L$GQ�{y�Q�w]uX[�IW�}�=r���˭$�'��Pi\�3i�ةԐS��Ú�?��)�Ń���`O�!�2�3��8�'�J�z2Wr:"��b�S53lɦ��~��	�3�;�D�Ix$L��1<��X�o����O8��ձ��N��%���Z�*�[J��e~��џD"�;����[���@iM\�T�Ż���o��bΒdXU2�T�ڝ�ˮZL�x�Jk�
��yWp�JG�������Wi��Z��|��@�eEp�\?v2��*)����r���:@�.�����Z_�BK/�b�\Q��� `�Wq1�q��2��k��:�ү�?K8���B�
�U��k��i\l�	��9V 9�q��P��S�U]&���8� 6��!kP���Ŷ<r��z��c�z[8?�$9v4��#��4��",'��ݝ��ڈ�����U��˵+�`��a�(ބ=	r�H�ȝ6�2E�]�].���(I��F�g_0��I�˘?Zq�{p�4������M�
Eu&y2
~xӻTt
T6��kU�8هQ	բnЊϷ؝z�[�T���;_�0�����@{꫑<��;&o�wUV�h7 �G�M0�Oã��I���O�+vN2�����͂���f���f�'���5M6u|�M���J靻3� �a4	:g.VPD�C��\�ߧ��Ե������^c��K�5Wfp��Y=	�ʖf��PH�c�D	�=�[�4!у,Gn�ẗ́���|�}N�Q�6�=�7��׀3���q9t~}���;I;����g��F{���r�" S��yg���p����ꙛðx��.�(5T��Z�)������5��-1f@�����n#gA�2æ���������]�;zq-�+Ww|�Cy�U��R�8�,�]�bQH=�W[H`���m;fƻ�:7���E�'����Y3M��Fq���P0$ut��՟G�Zb��_$�[e�FwXe~KK��Vv�]`f]�VM�����t�{1��J��SM�%��
�A���ɜ|��<
�\�0�=p���b%�C_�"õ�|7Ĥ�pN���<U�}�Xs8��� ��X�NS���D��d�`4��� �W�	�˕�%;/��i��2�'�TR��gs�+������3[R��Q3[�f��X������づ���"G ���c����=��]�܌��ؙٍ�B����a�Y�i��������|�j�uV�>L�A�b)�J-��
-4bbb����u�D��P~np5��vQ
0A��0b|������J`h�o�o��=L�4��gh*$��D��t1xȦFL�뿵$7u�y�Mͨъ`���/@Մ� AK����d�?3]FP�U`��k�A�ȩ4�Рҳ�湚c:FL�4M �A)$�O��(�&!���s��i ;��'��)*�[v����˸B)��{~5$>$��Z�qNi�x��`:���R� �D?��GR�] @i�o�F�mq噕2�s;��9 O��i��:�L̺.��\_vJP�\
f��W���Jl�O���eQ�8,�K&����^C�丂I�v����E{{C�o�s��B��%���2}�L�V��`�E�-�K�i1������d�j<AoI�bs�BG���z-��ߦq~L�j�b�B]���D@D=�6[⪯\��o���?^N�#�z�̾�.\Js���[q�x�܏����➆��"��Q���7ϡ#�rGAok�����'����'32yJ �g~p����<:̮��^�&�!��
��L���Z�!DRj�4ݔ�Ŵ~��dLp�?ݜ���8ޣ5|�J�ܾ^����P�;�혆�khh�Z����М2)ٺ��c���K�����뗘oh:p��̀�Y��7$_(�؛�+s�`�w�2y��14}���)�:��ÏK�$�q�Ǵ�+�1�^U�y��������vҠ䀐�j]�<xuڳ8��.��)���7�<�<e��9���ᅺ"!�]܇��QH�߷d��{�꣒�Ǥ/�^�$;G����⇶Gs��������]�a���W)=4�T���P�jW�4/��9}趨�M���7���Y7���.�\`����<������W���TS7�X��3��֮@1]},C�1�Ѕ8��'���N1#�2g�A�[�Q��s2��9�	�$�>Ƚ�o�I�"��/8��)J̄M��%�v�xuD]���
�}��*��M��FW��49�;�dJ�)7RQ�_b��p��uw��Mj���=�j�R���T�+k�V���9�p	� ��5��3�UԶ�?��L�W�4}@6'+�ۘ��n���5LGi6�o*���"6&�c�S
�Qϵ�T�N�;z���zV��� �m�4�b�h ��j�=>�/�$Ȍ��P��%�]�j����|)�U��-&�ӒH�%ѭB}RV�����J��G��<K���}�e�D��'sO�}1[~$U�_8q��D��U��Q�@ͦ�d8Lʕ$^���"�>�Nr�#gЅ��+gq�p�P���s�$|�u���U���s�B�і�[l��6�	X���*��j;F���-]vr�E_p��<�A�*r�K�U����%@��!k�nC�Ht��#�|%�DJF�F뤒��k�,��7̸�+0:�P�d���5l:�vx�g�Z���b��"�X�*���i���h�2�,�!I:�$`z��dZc��h�ڗ�8�N�1�"�YR��qS�ׅ���[b@��I���:�����)Nz�S�F�z�\AJA��
۝v^�@gT�	��?b�%��b��{﵄/ж�M�wѥ9���Ə�����s����19A*җ���LW
0��oCZh^�#8*�k��� �2x�c#؝��ٖ�d
i�����m�Qv�릗0�1%}�����P %�ć������ı�� �?c�g��NY�4�J�R�൏H�J�i��o�ͮ�{!���4C����Ɋ��c�ԗ�:���!�����Z�X���셄�=�F�m*�r��i�ԇџ�=><�^;�֯�Na���=�q5�PP��y�[xC�O�/Z|�����j�b��G�߯�q*w�%Ҏ��4�"q]X���S��S�L�8M+�ƢZv&Z���&���	2���Ȟ�򂵒����J�b:�'���<VkO���~���Y�8��
�ކ;4���ap���ݢ5�&��\���b\�؄��,��*��S+�u ��z9��ƚ{�ezF�@wU�7�?G�2oa�\�}!pp�7���#)�O(��jwAI��ʼT?%j;<��zQ9"j:uġ;(,U�X���"�l`]қ�,S�g�~��F���W�ҳ�H^�LBt����E"�\~�A$�4�uϓA� �I��O���	���@ۥ�%��*m,;�H�}�Zj��oV��~C>�X�'�Z]-�^v�JE?D�S���o�2�ӂ��.P^�����t������o}���B��<d�x6��G�@�a��f(ת�:��cC�f=B^��Z��2���6����P��&K�����/34;]��{Ȃ��3��j!6^\�Z�~W�z�ޑ�[U����u{���ʺ|�3Ȉr�CG�'�����r�c1R�u�����ZZ �!bge�ZX����
��p9GJ�t$p�PZF@I�~4n<��,*�l��5WOH���<X�X2f[�����ht#z�*<��UB0�h]�<."����An̔��$>�����]T��hJ���ߦ�FuYh�|���Ԍ0`���%��t�) �e�`���_4*
� �Y���7_�Q�{��|EtE
��������.�#�QtlL28wZ�)�Ï��sv�(SW>3�m��$�c[0S!�u�d�C�Sl�Kl��{m���o9�~����*
�k��L~Xʽ����4r���G��������o�43���Q���툿��1���(�Ls�S"��w�u԰�)Ӿ�+�_��E���Tp�A���r�bX�D��P,@x�bȖ/���vR@��̭��'듐���E�]2�D��ϵ���#	t~,��I���8�ݥh4� qQ�ޏQD3��_2������*ټO�����F�/�
�&!��́jM#�7���B���^�"T��%bzR�����~7��� �T4�%'���>w`������ի&��b/^6m'U��uMq
��[<,N-����F�4�@zǂqK$��=}��GF��y�{�2�;�]�vh	 �8��P�΂2n�f/�-��0F����8
��X��MR@������� ��]��aP���q�(c�-v��-�馗+����LZ�W�Va�O�u���&��. @|�����H�����3+�w	��F���j?5Nr_j�wv` �`%$�jj⩓F�!�f�<Toԃtڑi}�/�a�6į�yӭfO��\V��{P�k#���HJ&l_���gX�����z�v�2�!�V�R��X�����񥥁f�	`*�4�<�3��w��f��%>���ɣa5ī'�����Դ����)A��xA���I.v4�m	�dE���>w6(���1$�ѧk� 	Tmk��k�K���Q\j��e��8�jϳӑ����s]����0��q��]�T\	��:�����HV��0�&��.hҧ}��Fؖk�l�.or�w����J���{S��l��ila؃����:�Q�
Bdq�(/r���\���O`�?x O��Nmyl�
	�1끘�H��-�^F	�%u��h��@��>UQR�1R3s�~��V�i�B�IXf��.�~���ω���!�KΗ?=��YoE�d�g'���?���H�5�]2�b� �<-JB)Xԭ���ǘ���6��E|y��.�*�M����?'*kD<��.z��zn�#Vw�-_�C5_Q,㜍����D�i�����-�2�	�n���ȍ�B��7��D�X�ߤN\�h�O��
,]t0>C���uO�����[�F���v4xw��8o/�FU�ƖA��"�
l/���
��'��d�d#�L�<���xZ)u�?�g]��b
H����2�fN�:��/��^s�ʳ��E��Nhw��3oƮE0̿b�c��Y�9^��ŷ�֘��#3�q�L .������0�3ʾ�@q{4�$K�ݧe��$��Nb4����WPr�&BͰ3�H�+�:����)!uk�����j��=��V䰦��G�x�1 v5
��~�Pp�c�%v�~]��?-M�Y�805oBc7b�h�6p�̇���`�,�7���r޳6yy+�o?|�ݤ��b'�v0�Um�0�GCo��ڛ/2�e�L�&{\�L�7�1v�@��6ŗ�Œ�4���ֻ�9^H}���4)B�#hEZ�b��a���e�j	�ԛe\�WM�n��rѴe첇"1�JdF\(�Y��I�fr�w�|	R�S�͓��Æ� ���Z_�4�.��?�6�|�JK��KV�j�&��sEn�O7��Ă������p13 ��.6�,k�O��׮d��0&�����Q�
��mt��c�zB��͏٨�b���	>�_T�1�@���T�yT�5�!@1��m�vL|���܀�	�3���x�A��TN�OU��GO���v�*0OʤC�RF�!�ze�'���(����,����ta�o��~�:���'����@
�R`�%��52DE�������y�`���+_Շ���y����.p[Qo`C���\E
]r��"[Uc�;���V�����@��]����M��7qL�t�_T7�9��&�p(� �b�uO6�_�;���s���P�a�������T��qc��y؎�(�2��0����ړ��!�ە�b��d(k1��@% !۬iD[(��S
CC �W��=|��{��q�S����d�z��<�2l�q��q��f�(�����E#s����QUD��,U����ґ����������Y�9y��̌�m���E��\�$��i�1�RSU���+���
�H�:�ޡȟF�-,�gb�Y����8i,.;Җ���ߛ�"�.9�!�>� �TH������iA��k��)RS<Ӱ{�#
���`��.��,��Ohl�$ͭ��FCJ����T�&���x�ߑ�-DZ�>:�>���y�<��]�:0�κFk�/�k�� `x5����s_a��P�5��ɰ���H��RdO��׽�ܠ�h7�AH���6[��!S7`,"/|���E�v�#�2�i@X=w�4=sUQ��7)�Rʭ����!�_�%���7�>'���d�d��"�2��>��t�M:A����l�ѽB������bNA�xb�kY���~��ԩ�P��
u��(Lh�f R�V�[Xntj5�G\
q��қ� KW�P���_�%�ʤ�r��r�x�Rw�3Vjڑ�{#����]��J:7������k��%E?��H���"�SҩTS�/��X�Yف��6��UV�S�PU���zF��.�z����G0q5�겼����7�^� vF��� ��'����T�	�1u���M�j���T�Q�#������)L���L�q ��F����D?I��\�E2���O�n@�ݬ"Ξ;d��a�Y��Z�h�K1Z%$���d�UFGb�I�X�F]ÔjʵmI�YC�Ž���u1���9�c�*��JU�I)ޅki��2�>!F�g� � Ʉ���4�h�NϪ1���q�݃�Z�揅e2OH+�1��f*��&��a*Uu�ձx����{�LDN��B+~8�������sD����-9�a� <�0߂��D
(F=�O�`~���y*��a�m �t�������W����Z�=�7G�{��>Ո=���ٽze�xS9d+H�HW4����J��Lݐ�M2���e;���ݖp�� ~���L����U$��Y�  �sf�M�������8�.����#��M[u�o���ض��|0ëm��㣸j4��rzd3��#w�~.q�G�ö%��`����8��Nˣ!�k!��X>��MYb�D���<~�J:�}p+O��Q�Aǿ8$�b�Rgg8kh@v��l}&�m��Uʁ�H%�h�vh�U%'͗}S������íI��������f������Y����3��1�RM)�fJ��� �a�½�_4��p5��ܶ���F��x?�N�h�	8�n����;�K�q�?b�}Z�q�)�+,���c�j�o�{��qX>t���K�y�j�'�g�R��H�>p��� ���h3*[�j��JV���G=|��+�p#�X��j.T��m���L�u,��y�ш�I^�<���e�} �~Mel��`�ܪDY9��G�4\ ��|��1�����@b��o��c�����ֶ�(7^U�¶S��Hv�Ha���N )��B��A���/�d�\>#r��D���k��ϟx��"�uYT�,���#E��:<�*���3|��TT"���P��_���">XCR%vˤ��~*�uT�lOYyk��2�*��o�|7���bX?`�1�\-FO��)��b.?�l�NB��e�����ٟ�M�#�g�hL@�˔J&���eN����MU�9�C��.� ��҃���]�Ұ�� �-�[���_��k൪�sf�噰ØN;�T��
��o��Tb3\���Ȳ ΀Y�s�Wbel�YP��'$8h�F-D֔G��b��Ԭ��$S�5��N[�K~w���X\ޟ�Y7��|�{��!I�����y��T�{��Nb���4�JAO�\�[�fF���l�ʴ�����l��s8�6��j���SF����gޥ��o�AJR5�8����TԘџl�i��W7Kս��$�X
���P�B�<���b�Ր*���g�T:��/��\��|f�%@A���~� �vf�D%�ʿ���}�ZG?�{N)�$���Cɱf-���B�&�[u�8�i��|C@���=8��-�����z�"�/�5w p�&eR%�ѣ�Rc�B zD���Ig�c�,�[5�m�8f����r���s^�,�!�������iɴz��/;�WA
� �m�*�Я\�/��`ĕHЛ�������m,u�����V�/pNb��/%���|hr��W/ޕ���)���h�����U�ڸ;3�7���53@,�T6ztF��Ӽ?tӤ\k���¡.Fp$�9��$�s��ü�%:�	������QgEӨt��a�����'Gl4U����+W�m�⍢O`��b�t+�$@̹�&��|��#��t�dG���mE%!;N�5u��W�A�{�]��e�>e���2"6"��*�2����n:㻯��5�o	0���kl�k��1^�A����� ��p�����)n�����f�ܲ	`x�2�J�k�`;c�y��uV�p��E�]5ɿ�悁,h��.:.�9C�K��*K�U1��M.ؐ��`:����`�����;�ӟ�f6=_�+З�����p����;FfJ*���_<�6MR�y����g�uXYLALM���z���p�5�X���̑Z�*O3�Q_���@�~۾�qZ���X�PM2Xլqn��������7����A�^����_�qZ��?OD1Q�+&��N�����U��i�����U�*��☾�i�k�^��R̯�Y� `DM�sS?;0���u:am���ג��ئ��n���>.����$5�X+�9Y� �pb�,�}��=~9B��񸄴�4��2�B�c���|��&%���b��+�������q�3�cE�����c�u3S���#��_��[O����ҨP��$� ^�פTh>�vN�.#\�!��+}�>��F�t�p�O�֪��0T�}�&�U0�\�AGh�#N����/�W�,�~�s՟�K��:�5Xj�vC��ǯ+$g�ʥ�Ө���P�s�Z����Z�?��ʏ�S�3e�ʮ�=c�D�I�7?�ܪ{#�HG��n�VB����CR� Ox�e���L�7y�*�9�9�R��0�:������	b%D��</��Oa/L���4>�5��TB�o�R��S8�� �"a7���Y��<`I��B�<�BeciU�@8���:��	������r�{�'Ӧn?�'�mON�ZEn��'1Xz 	&f�V���J���@�H�pA5,x�w���OS)� �Ԛ	a���e�g����0��g�/�2�)T��kga=y�����P�/
��~Ǿ�Kc�d6�U�����v_v��%LAL��Q�*F:���������(e��=�gK�@��m����
CE�wU_�����o	�Sk�1HG(�#��ܙs��j���ɫ�a�Ț�N�s%�
����A��q�m���%�s��TF����sU$9�FH2�x'�¾�LR`3�,�3|�X����#��C9��D��l2���%���7+�00��Ƽp���c��:��<9[��m��E��l�����������h{���F�,#��b'����z����<��.�7�OkWM��)˼Q.Ag���Oa�=7ᬻb����p���.���f\rH�d!w��
�W2�`ר�0��a�������W҄��˰����$D7jو\���cۀP��Md`Hv��G�!Dzך��f�x@���[�г�Ӷ>��t��*q�%e]p����h��3=���P���SD������x!'�w��Oi/��Ʀ�6�^<����t��ג�Z�������$v�$K9�����_CR�^+����U��ܻz`��ڀ�a��!Y�|d������ɨ�$o�a2�t��u�1�sJ�1#�*q��?�z�4�m�0{��S4�^�m�<��L�	ZT�9��L��@ۨ���f��8|LyTH�e�:�;�����WS�� ���SĠ�[�k�:˯���l<0�0��jܔ�T�_x��\����9W���F�Maq��E�C��ݥ��a�7`8E;�ڟ�S�-K��8�Q�\�4j�r���r2���g�d���l�Ջ,U4B1D�5�@�j�s�b>wb76@�rN���絥�̜ݚj�-5?^�"л��.X$�	�;��0�5��Z����V6�dG!uy�'[x��n��rՒA�g; ��&0�2��;� �4V����m�[x48�W�^���r���nT��-rl5L9U��̿b(��3?�4�y����H��P�3�`����T`�r���PT7�;�!����O�m�|ӣ���U��3r����s�����Ƥ��&���A�u5l�f2r�QU_HXv��9B��!r�����=�{�O�ܝV"l�Xi�S�E��Xr,��c|���p�,�C�	��}Z�"�}�UN��&
��h~��s}���(�`������1\o��0���cI*ڑ�ݥb���ig�[/����Qtke�)x�Y�I�8��ߚ�lh{�޸��8
ym1�F�Q���d;�a��r��)�{�ʂ`�'qԝ���e+Ɏ�@�^�fu����wl�T�*��"����ó��G4��ԲCe���?�=�ь���鈛�Zuڍ��{1K�(D`�6Ÿv�j�Ԅr��� ]V(b��=v�:^��R Q1���fz$ sKNx��D���S��N&�V�F%�%��*�U��G������ [�}e#}ȇ�N�D��Lш=_a��A�/a`�H�D�\� FJ��2B?ɢ���X�%�8υ�;)?~�]��o �v2��	 ���Zy�W���,a���� a�a3V�	���WºLS%A�DI�̾5L�c/�lS�����T	ߪ�x���g �{������n��O�z3G��s
�ue͂_)桉21��ˑrvgl�|�ˈ��TqpE����m��!�+� �,e��6+Ҷ�Hc,$n`0���Hj�+:���k���yc�#~o$�q�Z���1z�)kG�ϠI�����O☥�<��O,wN��:(�Xr���Ƚ�甁G��xnr�l�nIN��l;�o�¾n���SYm�/5�����]읷��b��L�#Ý�X�G��f,^K<��O]�uL���ﻊ��W 0V�l��4�$N[FJ�lZ���7��af�?�М˚�%�h�]�,�,-��;c�S���� ��U��}A�Vbac�J��93�7G�UP緎�eV�ߊ9#}5� ���j rpKN��Q �;��{���&O������Nqyؐ����&��`��6�������4��7O=�j���9�f8ئ���7�V�j�"��|�S
��rb}�>�8�I}[�Z�5�c��6���Pr��`e:rȁ6��[Ÿ�������q�3�`D'����,֛i��,��j�J\=�`"��#��x2��cZ_�Ø1�-�ދ3�M⁋��b�΀�u��p�e��>�������:7w�e��'0��cRDG>)Ȏ�}����x��:���K����5�l���Q8�?�}��eAX��O�S��d�j��m%|�qeo���w�XtC�����H��ழQW��H�Z}q�Z�kT�("6A�[���(<�F��`��+�A���)���W��,��-֑
���o̸�1��/����N�u;6�XR�|���c���3�u��Q�u�xr��K�qE�{O�������gA�P�q �p��=��c�bm��7��X���˽7�O3��[��9�#���0~�`.� $|��G�gZ�F^Ĺ��&��y�����י8�-=�d[�>��gA�*���o��ǒ&�������AN}�Z���w�OTo��R='�}�|�E�=�ZN5��_ �O��\K��&:n��[�������DAw^,q%v�M�;i<H���Oe��#�h�F�
��m�Y�dl����>r�t~��@!D��h���+w��sN[�{��)��?ю�nqT����#���15'Gr�`f����g%4��/#kå�
�6�Bn��8�Em͔.�ٔ�Òޱ��iG4]��������So7�/r�~'D |QΥ"�|��ܡ�K�v�-��Ta�\6�u#kam�C�O�s��Ae1WnA�����i�U�J�φ¯R���3�q��]����YX||���T�&�o���}�ٸ���M��������@J���Έ�cw��P�͊�A]���RU%�[!՟��;�0wR��W-�>�#5L�~<A6��0����&����68r�k��*�D�0�P�1��]��p?T��Tv&1�<n̎)��*
�Ĕ���#�U�����^3��M���v��5��}��Ö��o���У�.`~�]qA4}�m������#Ϸ�:��}�\�Nי)��C��t�����m�_���ضض�8%�H�^*�$3w��m����x-�R�������!�ݹ���<:�P����C�ssI���1Ѝe.*�fh��C�aNa��dx��B�,F$=Mƍ-�Wl4|���! ��lm�����k�c[���*E7���c+4BM�-�q��$�>�'����6l(.�[j��m�����3og�!�|-��&%P/i9ޘ�&VS�)ꕣ*�#�^���A*����9�x���."	�E��:R�������z�9N�	r��� �	�6��w^�7�c\�� H�_e�l�1� J4�GF�'����Z�|,�qX/�!R�z�z�eC>v���׳�tj(A�B]ؽ�٬MX5���Z�jR��S٥���n��4�Z�)�r#\��6<�����\��ρ��ӥ�C�i�ОEۮ����"�Y����o|泿��E|Խ�Bd��_�f������F!9���]֢�n���w	V\��9Q �;SdH�8*H���u<�~5�&R&!�_�"<�]���O���t���q�w�p�|�M���o3
���FK�V`ժx�d0�,x]������>83�KV��4�E�˝��������-�X��7�b$߼{�%���BB�X䰟�go1�G����gG���� G5	J� L���JL�f�D���n�'��K~�L�2v�v�̐)��y���Ƀ��R%�f�E'~� +����7A?bt��N}U��`���݄��Ȥ^jO�Z\����j͛��l��n��>I%;����ؤ��)�]k�]pJ�ϖ�[�tQ�Z,'�D�PA�9.�h���ie1D��)`V����6�*��{�@��[T�Ǐ�il� �b�CG0�#r���_��_΃xC�pݫ���DkـpBގay�ǄI�!,�xzhI��.�T�C:�y0R�!����j���߈Ը�^n�w��܍_��D���"E8SS�"��>`�`�qij�sv�҈FR4t(W_�B�^��;c�Fm��TRگ�2���J�*X+��7j#sf�ow�H<��z�p*��0��F���0�a3"{�T�90�F�����x�����0r�΍t$�p�����)Bn~�����<�
�-��c�Rk�tǶ/���J�� ;�e'���i�́�t���F��Pܹ�m���������s����L�Yr��W�j� `&S����Х�6����'}?e y���P�c<^�2Pp�,��ܯ_��V��gY�#k'���	��pSq��Z���tT�K?�Mv̉�5R Ւ}0BfK�=��G���e�p����[��G�P���vvo���\��z��[������K��.z��k��\��1h4�Tr��e��"JímnCk�'�y��?�u��Lۀ�:"��w�.|v>�T�N�"�l�y�^�_�TJD�s�2nf8E����ț-T@f~�_>o�	�6K��U"8��$g8�v靇ji�%�Qg����&��Q�RdV��$������=^����|�Z3o3e�A[��p��e��iU���܄S6��lOk��^�W>V9PgG�����b6����CR���i��{��z5�����|E��,>�=f9���"Jm��]�:�^� ?1GO�O��Z�H���^��Ҭ����L�i��+��1���)W<� C*LW{#E�@��u�@'�0 IV��'����;�fT�[�|��IԒu�͵�JQ�k�V�nlM�H=�\}�4t,S��rh7�d���Y��  �ȟQSѯM�����[�Pr�-w�9Mm]
#�J��Fܚ���s�`�� 8_m�r�,P��8�H�5s ��
>c5��Ũ��sr\m;[ǘ1�Hr9��n�_��|��	L�a00��>{���s��Slv��WͻX���M:���nE&~|l���G9,#�qk.�s3����b�%l�{8����e�7Op���V R�\>	�Qwq������xʟB�����\]��ȍq/��rt)���1���IS+��D�m�D�D�^4ߔ}�Fql�ƍ&��d�
���yV� }���%�A9��2w�G�����F�(k��$P�ܵ�Ϳ&ky~�J��6�HMK�+ܽ� �.EO�6�$��0s�v��� �+>v��,F�|b�.`��K~Y��a�)Z|<5��]>�k�{��gY�s�I`�~q2��Ŭʦ�E�Z:���W�p��@;�>`��[�����K�5yI�p���W��iQyGqGMM�G-��0O ���L����uvf�R��g5ZZ��H�ᙽ!��D�6�I���tx��욾�m���$�9t�^y���$u����5&�<��ua��@��)E���F`Ӫ�<vM�9@n<l��ix3Y���(d���9����M�F7P��
 �ӥ�1�B=}]����9��k\�Y�W���n}���+��L"���s]p+H:��0s�w��W�U�Q˓XDk���L�vLi����f8�,���ۅ��6�Õ�n��1�K�E1��[еY����x=R�u�]�/����mX�я�1��qv���r s]�v�i
;�p�V(���9����>M������B;��C�R!��3l!�E�p�����_:5o_dd�!�v�f����i�I'͔J.,��w�S[������=����t��Zk��z�//��OSq굲3GM����J���w#0d@q��e�﵂v���;Z)���a�K\�è� 4<ˋM�-pF��NG�|���xE���^V�r�;ߐ��qBNw|�'��~";�`�kP�ȷ�d{��{�~LU���謭�9���1�`�
�y�t��aS�����z�]'ڗS�v��"v��f������wZ���	�?���(� v�7M�E��t45�;A(��DI��4I@7A^WͅO�Q�n��u.=B�I
Н�w3i���-��s��_��6�&axb�����=�׆5{T#�g#��:�H�r��9�׻�+ꄕqt�u1�}��O�&��DR��@��ك�8�\�Eoo���i'�q$���l_ֲ�]�*F>oZ�
�P{��I\b�v�I����+ρ|8��6� �l;���g�k�F'@�j1�W�H�eAFP��,�~5YΩߏRl� �DH
���=�OT��!������3��b]e����j��0���#��wQ�S�z�P E���K���f7_������#Y��,��W%u�nN��Y��#�������ҝr%C�|:L�?w���?�5�ћ�4
�W��A=;���Q�Zv���z_'X`���FP�vC@�|W�⡹�o�M��n{��㒪�Vb;b��\�	����dAf��l���a�p�K�v�r��2�a`�+'���4l�sԮ��p��T�~U5
�}�I��E�P�$!k_1R��nW�L�bN��w����	�v�]���z'}[ؽb����%�e���k�D4���|m'��<�@�ؒ\װ2;�3��U�6�J�p�W����w�r,Ѿ�\�����AE�&<&�pSHA�Fb���m��I�o�M��큽�ɖWˈ[���xl
+�:5��L6HZ��s���>l�e�Q�W�|���f�_���鄩�\�c��f�r}�{��"bG\өø���4314H^���Ӣ)�y[�bL������{DdB�����2*f��9>�J����Kh1�(/�-����T�%��N�6���+�,����M�����UO?�e�v�9^����
VU9�"Hy�n��؊M�|$N������6aw�sf~�ϻ[م���>��Sѯj�9q�,$��e�MA2(�4��:W ����0�o�dV����ܷj]С��K�:e�tc� �����<'�Qg����gH���{r����N臃1;�	����?b��5��t�9�	��Ms��`���h �5��o��ϯ(�7Y�ŷǢ�aҭ�b���.G��7o����J.�[9�	���n�fM�����]9��<ײe��ɠ&�1yr���9ے�I_=��,h�/�L&�������s}G�������/�����q�Q��72,��N�:�Q�;�B��e�~�On�`��E�봦l>w�a�;�i^P�A�'�������|�>}%�n�JH�2��c)�Cg�XJfB����H����}w��h����(|x"�d�?�nLN+�&
D�*��j;�l�;.}�2^R�����?E���s:�u=�,+�Ӧ�u��Y��I(��p��Q�Urd/�j��z'r��х�S��k}+G��<���*�m%3��ݼ�gf�i���7Kq��E�]'@�α}��*��ܜ���=�8��w������Ў?��2ϰ�.��݊�.u@��:]�I��V�:q��-��ح�;c�'��!-D�%;�.&.��*&8^����H�V��s(��*��g�ٷv���iӡ�)�~4b���0��l3�)`�R�7X�%哬M��v�[�V؛��HUy���T7,�Y��ć�aW")g���z�˱b�?X¢�`�tp��ր�����Yeo���HP��Uc�K�4�P'�ڍ�'
�i�M[lH��z�7��_B���m���Z�����=��q���>�_�!�����E�y��;��o��-i��hf��y�W�A}x��E]),���.��}����K���=�z5����|��p'|�����b���#[��� ����ڕd{�V}"���MwT���}D�j�ly��H��,�G��#z��c{�d���,Q�D `���RP�]̈́JZ���o��vX�>ğaҿ�k.��Po³R⣍���Wd%4 ������d������ڜC���V��J�"��/�f/�_�C�`�?�C����	cT���6]M�柙�Jc��0Y��2�_�v�F#��8�rAnVU"N��:�-TM��o���|!9{s@[�/��� ��^�`!#��b,x0��B�/����jxBU����"��n�ɂ�ms𘏲R�����_}�Cq��3)�%���T�Lq�n.n����a���2E0*{�.�DR�TD����c���dقߖ�0�6&\p�7au}u%;	�	"6�J���MaC�{��$�IB	���1�w��;)���j�&'��H�Z�R��H9Q�?~1f��R�E~�~��}BD���җ� �j�)�pP���d�-tH��oӺ���V
	��^5�KX}�[�8Pjl�Zs΀#V/$�b���\�U��r�X>Tϼ)���0:	�^���xJ۟Hxxj���2�_N�˾Cya11sH'VՠT/lw�B����f�1��9:&ig�E9�~�ʫ�e"徯���%�d�"����������9<y�fz�"��
�*[�����1�闉?��5ΰ�@$X�;��(ϱv�n2�B�&zܶ�y'�����zM\�uu��Bq����6����RQ�6��8��+�l|��+]�U�h�A캔�w�ǣh��/��4�||Q?a{��^�Σp6{&�ǹ��8�R2�_a��"��x|@,���
�Da[:pފH������a&z���]�i�'ט�`t`����
L��<��u��ko�qfR�F����i����bY���6�Kj�s¯��m��Wߒ������q�EC�VP��OYL�~ݟ>�1K��N�-G�9[�[��4	�_��ʨo6�c�-;��c�aiynh�j&�KU��p��Y�+6	��x��P�H��zFGo��࣯�a��q�� C̳��,.WӸ\����T��ڠ�`���Í��[	�i?�荵��vcIb������7/��6#�b�b�$�k����S��qn�|"�3�a���wn	M	D���9Yl��QL ܀�Pc���Qoe|��Q�}n�,�����玂sD���m�Z�,nܺ"h6���L���	l{�ꌿ6��^�w[�������r��K�1^M�q~^a����Ǯ�M�K���t���_p�60k�pnZѬ3�y�'q��]���(.ʛ8}��=L�
�urA�iG޷z��Y��K�N9�!��X���ѩ4@=��c\NcRμtS����ú5d:� vI��������P��"D�L���^&��`U`��}3y3�ЕN6�(ٵ�?�����qZb�ӣ�� �و=<�$�> ���c�\�ֿ:k�����}Ǎu/oo�
�T�
l�7g76�X�#�����D�������׬{n����.0<�"O\�KE�ƫ����^4�_�	M�lMΜ[y���fc��k���.�7�ߥFx��HH��S��A�~2��岐��V}Pm�i88��Wq ��ѯ�d�T6�EW`��\\9�\'�n�����vM�g�
A�B�T������P����4�N1�L�lC�� T$������Ã���z����X�U�E�/��	�x�m�
�j֥�� �dLok}^{���h���%�U�U�a&�߱{�NG���f�V�Ns��Ӫ�-��jR;�O �Ob���[��7Ȣl��(7Qi+rr�����檞<�K\���� Q�2�� Y#��S���[C�:�d�#�a�]7���W������F$�B�гw�`��a~�[)���~t�(>�k%��ce[��N
<	������qk�쇆A�<�t/���c7]��}K;�d7�.u�O����Yb���r����i�Gߖ�x����q'��!����RS (��
 �7���.&�Jb'Ƭ;��_�1�♄�ΠԀO�J�k�G���qZ#�g��U���
�# �.�Lڏ���I�b��M=(_J����3��	��m��eKң_@�o���܄�Bn�w|�uM�0��Ρ��)0a�xQ`Y�3�i�"~i��W�7�y�Y���跱������k���;��O��c�3�6��`��F������2�/��q�����6��9���;؉�4��{���4#b���7��K1�����-b�w��xL����X{���l����xE���u�R!�,�p3 �'��8�h����)�/piEP�Y�f!��2��c�|�1� U��Z �0�'�6������l�{:���h�\Re�tY�]����J벼�z�|m|����AI5[���Z�,���5#(����ٻx���oӥdB�wW7�S
�8j��r�:v*|��;G���2)��Wr0h�sQֺ����Ot0<HM�
xW�㜙���-Ӛ��{%��&�5i2dm�&�Z��)	��Hf	�z�Rj���|��=�uV6=z4u䓈�YGF������G�'	M���Y�aҳ�'(���h�Ψ<��9��5��;�E�P�(���
o��#nK�������ծ�&Y�4uvj[�e����h��j�� r�NBIy���d(�p�g>���h�i��s44���ؾy�zx�e�@��q\|���o�e�`��D�s��)谩���S������}���ܔO�q#c8"c�q�Z��bȽ�կj�6��\�^=s�Ү�'kA�cRCT�<������PE��I�#��U�hlB4"ݾ��x�L9m\5���]W���b�(��#�_I�Y������0�Ӝ�~,�=m���X�!f�	��7:���H�pH�Gضna�	U�g�̽Hs�G�9�"����]�����btQ1��3(uA�u��q��^��-���Xi`�3.����7�盼��u���#�o����CL@�(�Dy���0{u��
y}��FM�1�[$���?���_.U�#�v��:m�jsvH�z���;N�A,=���c뻰�Pq����Tl�� �q�6�	�Y�;&�cg�z'�_�q���ʴ&� )^fC�`��P�����~R+�ɖ�!7TvFq��9��OT@0�����\-Ԭ���"����;y�~�{B<2p�0{��\歅�n��IO܇lK,Ҫ}|�t2��*�#��hR�5>�r&���1�W�%���C,�֑����/������T�[e[K�"1���0U4��S(�a I8�h1��ܚF˲ \(�
����d�.�I"
X1��� ye�M�d�i�E��B��<��qd[� ��?���0�2��qDxF������2Ǽ��K��=/ґ/3S��0�΀пh:�� j3�l����\���h8=����(�N=�����G�t���O�����7�%z\�]���_�,��L$*����ag��̲�q��E�);N��f�o�O�� i+2���[$�#�b=�A h�1�W�"�g*ր-UV�(�Fu�{��bn8�_&$����*�?�����3fv�8^g�L˺x�����^LB�hͮ������me�wY��J�J�ȨSyX�Z)��(�ɬ�A���m������$9a��"�����Th�/.�M�g�Q��:3lG<��C�Ĺ�p��έ���p����B��5|M�"�e/Q����hkD9�����%�0:�k�ÿ���x�5 ����n�z�y�y�4�T����"(�
X����ċ��U����h+N�;'���D�K!vg�[)g>B̲Ł�ck�)Bת���)ߊ��]�(��.�B��Qvx�#�C�7�1
$1S{�@���?�׸�N8o�.�zWb{c쐭cw��	��۝uG�!�{�����E#N�f�P��:Ћ�q)1�k�~��Q��ڙA�7|7z0��t���s��/�/7�c�hRT�+�>G�ʊEa �G��zw�-8����b�kb���,h5�N�^��mr]U��SI'�$��x��"r�m{�T�Hhs��L&�y��^Iz�<f���[�?մ<R��PQ5+��d� �I(]!�p$�M���	�۠h�᱕���_|y\�AZ�W�+�[���[���Φج���z�ͨ"o#�'�(�He�"���u�>+�34�~v"�8]��癨��g����i͋ec\��fv�_�2�*u s��%� �����e�.�:X�c��a�|���U�6����/|Ht/��{��j=�B�.��*���G��Kvn��
����QY-`�jӼD.)GgE����"�~��pFxh���芮��ȲaD�JNn�RU�L�ш��iW��R�NO�R��5
�u	�%�Z�rw�h����:g��U�Ac[�<?��~��I|�!�Œ�N���9�����%{�n߭�Q�Ń	Z7KJ���) ��fT�����Y�Z��\���o ��\��,ߍ����{콉���I����1��!fJ]Y�#0�֮^�����!qk0r�d0.�̀-Z�׹�z>·!ŻHY@-�F��/�`	�f�)C�r��{f�q�.�g�\�T5���ϸ��}M��F��K�1�>,�4��I���u�e2�|�
%��V㕳pgW���>�
#~�i <��㎡����H�>)|��`�H��Zv��80�X$�j�?�Lm<�&���B��<�L���/c|���I�O����N��*��r�4�5KH�j��w���
_W��&p0F�k��Bk^��A'��~((Ɲ��p��#�!���"]Լ�f�6��:����z�;(U�.��h���+���8A��my��
�|'�.�.�,�b��cu��G��ɉ��|HN�e����K9�lh��\���7�S��%*8�����W:��fr_��)���3�Z�g�t�ƈp�sy"k�;�kB|��Qur-!O,-������!�X�Pq��.�4�Ȣ�
�5�"���+u�N���Os0oM�. �1�&��s�ڹ�S FP�5�n���s�P�����3;�� ��?���gv��7J���ɺUf5�7�7K{wS�!�j� |��8b�FU4���K�B>�i�.0J��&��~��R���_x�B�~�ZT_�<TD�s��72��$�'}�$�7�
�pj�
,<+P�EA��1��kW����!0N�S��L3����2Bz�J�1����T"1�� �[�lJ��8��cr���R��:$J���V�g�����;m~0���1�4NWm�52ڤj9���2L�%�*�S���?�#I#��
�i`�KB�A����h��v]!�3Ź���zm�&�
^�>i7����Q��W:eb�(s�=�K=l���VȺ?��>�H�N٩(�9��i��p>����ʃ�ʖ-{�W)P?{ƈ �u Kꇠ��~�+]&�i��'j��y�'����K��쵌�r���T�2��IrQ�:c�Y��sV���΍���ξ�V&;MN��kA������L\���Ye�.�xh(���GJy�1=7���f(�г���]�ףfJ�Z�q���@��}�B�2M���F�>-�<��'H�ӕu}��$"/NR��O��'��G��lu�� ������Zw��{L�������I�C��Ґ��lH��T�>�]*-�V���7Bw�b�R� �;>��>��78y��Hd��P��y�fg��A���>6ʔ�2�:��;܍�R���&2͢�ju��AS��h<�?���|�SLK|&}$@ǋ.ښ���4�QC�i �; f\��8�O����i���nѡ�vK��D�֏�r'@����q�d���U�~l���7:�c٤K�����M��B����R���x�Pm|�@���W��]5�z��,>�Zѿ��K��}lX�Ƿ}g����b�'��vZ+��8����	s�j�8JL�:��i/C�Ƶ��ˣ�������G�ə�cr���һ�h�Y�V(U�I�~�<�z���uj;y�`�JW�g*�W�a0�����Z;�g�k�v"2UP��p�;8Q�Ϯy]ǻ,�*Z��
\��(�c��<��!m_��Ĉ��^��hb��&��
�c� )U�0�h��C+�o�����ʤ"�xR��z�`Y1"�H��$�p�a�l���T̠�iaFO[���r�n/e2u�yݣ>��g��0R ��'��[&��q���'ɑRP��Ə����Z�_fx>��N�C]�~��|��0�*��s�+E��4"�l-4�]���W��h�-���	H�3�&*>�'����U��[����?�֙m�H ��|]��M}��7�Uv<�_���38��L�-L�p��Ɠu�(D �sc�=渄Sw|�
f5ov�����t�/F��6 B�s垥Whw!ƚ���K5��(�.��VA�>�@S�CUƀ�5��||iYKX�[�V����ّoU�)�����E<6Ӈ�D��\B��اC�p,�)�}�}=��B8P��23R�j�n�)�_��0�^�s_L�VN_g4EFa���^�+�S�Z�	͊��+���%�#�rx�>Ne����%��_<�;Z� y�f�Q�3�&}����8Ա�F��0�?����Π�:3-'�w���Ms�Bi�8���9�_��g 7�@�\�Ɛo������\�u[�͞3Vڮ�Ok;���܌UO��'�R�@Xx��"��C����?&���T4�>�64(��KC���L�i��A�c��"�mPr����Mn�B������X���O*���AD������׹4���^׎�t{�_)f���c~���7bjx�#VN�"����*H�LlpY�'>端x����?�κE-����J��w��g��L��+� <�1�"i�̚�㱀��a[D��_�\I-e�p<Nko��W׾���ur�������������i3������_�A>>|�s�#�=��ps�����@h?����_à�,e+Р~��L�0��K�O~�ɸ��	���75��K��!� �"_끉�Gi7�<H	��.!��w]�9�RY@ꊃ@c_xų)�D�l5J �>%�71j�\������ }Q3��i/����Z3m�t���J��"�aE�����K��gs��%s���l�o���B��U-�Q���έ��qe�O���u����×:B ��K5l���U�-�٭�u�j�7��o��a,T���u�U���Փ:���mj��8���E��7�Y��3u�T���^ �����*�G� 0�SF�J4[���d#$Y�����͆猑� :�ZH���6�7��K�η�����\�P�~*w����]��:�u��gJ�T���Hx��"L^G���Er�{�6�t]����IQ��A�90��B�� �sZ)i���	5/Xy�u�����Ν�eVj��葉�1?Q0-��(�$����8�����*^�q
�<���a��Ch�#�Q��L�;6Y1J
�B^K�0,��Yw��G/����k7Ͽ�ؗc�����ua78�;hlۃC�3�+�˷�ӳ����M�:$�Ί��[΢�A@��	�E�&��S�4��&�늾��l��^��m����v�n<3��tEl��b��$W�!*��&ޥl�T�K�L�a�����!-�p�9�L�-,ɩRމ�U�w䧯pf�ݷ�Ï�t��!�"BO.�8L�_�u&�R�%�f��J�`��B��wy�a��<n(�Ɍ�ĭP��2*�I�O���:���@�2c����SK��ҽW;���Y�a�����E�\�Z��}��I�0������͋7S���N�1}b��iDeͪ֕Q����]w�q.IPYdm<���wSl����h���S9x���.I����@�:��w�3���۬0�&�E�d�U�VN
�7�KBS�J\��t(�Mh]G��R���]a!�Ҩ:^D�˂&"3�7���d��-�3�xF�$�D��&��{k�j�ʑ��!�.~��Rfu)�ax��
X��9�(U'F�o^��z(��o��G˕�M!�0?��薛!K�cX��ݎx���MNh����b�;��<�x��|�s�)& ((��%��)!j����1ɳ�)��~�jwO��]�M�d!�J���� �,�悀�j��1�?����7����X�KI��+��F��+!`5�z���1`�͹�%���'_���_u��b����_�N��[Oh�9�Qသ���؛$x[���'�U�\�?2Ic/��R�p��;aLzi��}�ۈ
<�V�P�I����V��Z݀���N�z�%����$J����W;��(���ڥ��"�z^�y3�XqQ5�Z�6���o(�*@����
q�.F�Exu����Z�v2V��!���u�sY��
��J�S$:X=0�;p���.*���eӠ����=u���j�& ��*��%�kΩ�lů}�xL���F���y�`8L�=�� �K/��z�lj�~|������VG}j��A�r���0�R�	���� d�hJ6<?�7���f�(�i��Ę�P&
�d�ќ�*\�� �*�,���/��p�����I�Oh��%��.q�/^�I�J��⚂�s��.!��"�G�I� �ڋ� �$y���V��Z�v�U��4�J**������B"����-<d���SN��Y���S�Cw�`���3��<��*N���׬���=>�3ב%�}��L`�k�\�>
x��W.F�J�'�<�N04�l*��bڄ�:�iR�����4͌�+x��LL&��)�[���7!Zu���i���0�B��=�P�Z#�懑�QOpU��]�t�Tp���.a]���Zïь�y����1�/��-_�24E�n
ee�qx'���f����ws��g����S,��[]#l<� �_�˵��A='G���ϏN�4�Pb��>Y4@��߆�5#�0Ԋ�u����r�0C�q�����}���Pܵ�El`��2���� ���5!����f��j/�U
��jNS��R~�~Z.�cC{��W��F�=�X�bT�ӝ�%G�s)�<\��15���h��r�Y=C�_L�s�P#�t�R�ql�"(q���#b�*���"ś=M^E@��"�Tn��lZM5	S�d�=�r��6�&x��E��s)����wȺ�Ò2O��o�zU��D_�(cD���/�/���pd�w�v�Z#KHR��+�z������I��V��toΔ�L�G����x�N�g��*Jt�k
�i�(�>Xv�)5�{ҝ|�IVlU�=���Q��b�&�:��h����L�z�����n�߿!�K���<|g3HZ��L4 �Z*���\���HW7�.L�f2F���ff MIV�Tڂ��,�Z����ʜ,!�����������K�^�R�-*ô� ����-���QrPF�H�ay�ހ��³Y������P/�囜���<B���ChP:;��<.��n�J?�%L�ն����L$p�;�PnG7�s!�}�k6��P���$����}B7�y|��K��/�e�J��>����o�[�hki������V֚�h������~��͸������y���n�S�C��})�h*���6���_Z����dB��
~��b��ha��kYA��п<�?�ݢLy�k��q�{ w����L�Xj��\�� s�l3�3%�O�	��ۧ�9�.i��~��F*�
3�hJ�;8��N!��D�����̶M�L��QiT��l#NQd���J�;�5�)>�Բ��>��H�L��0�`R�Sܩ���3Ȇ�M��Ev9h������(�	�^~���$Z�ܴq� UP��|���*��_"�c�G��;x]8u����L&>������e����k.=�vA;�MlycZE���<�x�	��v�V�ybщ"b�J~����/+�G`��SsI@���i�͎Q��`ְк�1�ǆ��C-D�X�`RK+��nEh��U�9�	w�7�k��'+�,�mץ��&�y� ��>s��?�cr��̷�YJ�.�>�v�fԛ��@��6�ӎy��|\�{Tق������R���,#�c&Ä��G�r�y{��\}+��rbn �
˔��u�%���[ީ�+!�9饦r*�T#��$Ù"z4���[�M��΅���:���[�c�r��埸�hW��?C��"�~���j����$��_�q��3��w�����,�<����s�� �e9»�^À�V�-Ĵ\͘Q�4�n�$���A�2�N[�=�e=m<ήq���Ǖ[�L�">3��hkH�g.Y�[�ʠ~,E �A�f��_-���3a�?M
l1Q��ŀnB�m(HRŅ�����"�8��yf�P�A	]�
��q�*j�������TG��QI�F_�1������R�O&y�����[��d��� CdL��e�����l���rjAE�6R^����>$�D/>�ԎiŒ87��E�``;_�c�@�QZ��nJ0�_
�yu� V��2Z]A!���u�[y�l[��)��/��%����/��~��T�>/�B�{|妩��ZP�h�ȿ�,��k���H(�����
YBx?�)�_����2��	E(�f ��w�ZxڜV8oQ#��3qp�� 2�h�^�W-�~�볇��Pg:���ޡ�I�g�Z���W�e���m8�+����w�B�_�[j:��48�YNfh���G���b�����ڝ�0�mʊ��G��2���</�]�2X'R�WH���a&��6�0QQ�2�W���t�uu��Dw ��ـ��&�����G�w�ǜ�����K���-�
5�}	;�Vq�����綱L���䣣��+p��I��_����b�*5���<3'uZ��Q-�g6UueM[֦:5�b͡'S���N�R����- ��\y�v����m��D��YG���v�p9��&��a$&�yr�V�U�.ި^#M(��	�c-�Ƀ(��?�A���^T5��~�Do�������U��[/��ZͺhAɫ%EpAH|P
j����07�.0�����pH��x?4�y8��_�n=ǭ̓�z�Y0��3��T�H+/��[�.��bOў�-��iD����q�	����1�G�+CX0T�v|��#^ܕ�VhC�<�dO��^��8H	`�*|������)Lt�2H�r2���iF�Y�0J�Ċ��NY�� 	��{�U�`�]��g�p��-�*5Ǒ�8�G��`�:�ॗF��?�!.@*�ޱws �Xyx��O)�L��I�kw!&��c��J�z����i^E}_����_j���7�N��@��OUX�~oX��|)�<�tmSg�|��4�y����u�
d ���_,k�t�����݅c�i�q������Px����t5�&�=���N�����k�O|��#K���Ⲱ6�3kH���f��Q�)d��El�H�ᗔ���"`�
2IC�)��
!�O-����_��S+�W�`Ս9vODYai�>ۓ9Iܼ!��l:�/Xqj�kՅ�ܙ*j�P����Y��K�iRZ������YM��y':�i�ށ0#&����nw?C��d�th��Rg��� Q�S��_�NG�F>\X[$a2E��`3�g9�1���I�a3M����>�a���a�������|U3�Vm��m�m���(C�Ԏ��	�>R{�� +�&anө�CShͿv��H��_�ű�����v���䗪rE�fuh��N|5mɼ��vs#�����������}>Q �eլ�+$ �P@F���/��#��jM��߳�6��`��s5�y���^A���ba��fk�v8��ĉ&0���`9�L�U8�m��5y�h��3����a5�� �%7[MQה��=G2�p�gr�$���E�A��諟B���E��h�1N�&_���zAǼ�=���3����1Qfu 4���Zg��ƣE�5�AFTs����M���#ޗF�-#K�b��⾚c�a�������\�W��3��}�b��wl�	W*���c��SϪ���	q1��r��@�����:�L�0�˗A��\ot�[��U��cH�ā�-6��. f�;��2����D���-#�y�4�m��$Gm�Tj�I���`vM!`\q��{�ϤDh�/C��fMf��d���b���<-w6���ZR��<�����5���U������ʯ�6�Ă�P��=�\h��5�����D0��d�Z��&H#_�n�pIjz���k��%���[` '�r$�� F ��c��]��:(_�k����|�/���M��@bv�o��G"�4�V���v}�A����F���f��/d�ު_�\0Tj#~�K��(Hk��Y}��ɝ�I�jX�.֘��ר�e ��mg��<�]i1����kq�'�<�i�S�vi�6F��aˋW2�]���_�A�aX%v��9T�qJ�%��	e�>VF ��Ϻ��
�HQ�;P��~j�C�[t~)�Γ��(LY "<2��3�� �c}_3A�Jf�t��2�pgv�7FzG��qY���m�_���U���,�d���5p"�&����A@(q��91c����=j���M�#���h�W�P��	i��"��.�q0nf�Y� ����
���lmN��;Qs���Y���i�_��W���c�ji
���sI�Y���Dw�Ppv.I)9W3��@u�ˊ��u� �	��:�W������2κ�a��~�u��X��	�jYa?���5�ŵ����Τ;'�������g�WV�`#��Y��e��N��Y��s�!��%���u��=�>�?���d�	�e�ɾJ�訚D����� ݎ��@mğ�Vp��w#a��;��jj`N���_����fڤ�Ah�sʇ��㲃�vJ���b�#�k?9��V���9 �D����#dg�am��Z :�r��fH��`:�Y)�f�t�'����S��p\/�k����WyۥK8NX���*R'hW���>��clճ嘃��%��K��J �E�dV�:�B�R�p B��u�	(�T����M�:G[��G�͕��K%%��G�8	�����e�������[��U��)�����nb�w�R[4�82R
�.|�h��#��*��.,�e7�^�/w�����y��Fڭ�ـOAlK���1P�v�����(���t �BLo��h	�PI�����*�a�>x�$��� f�٨Qu��y����H ���ǘ����U�Zn쿔��JI���u�RI�ϊ.p��ɬ S��q�j׉��ӵ�
��$��P�mY�����bsهp��T«8��Z�Cd�w׭��P8f���>����s�`�X$4������Y�#��������ע�^��%d�"`d��J�|��I��^�{�diLk�:����ܶ0* L]�m86r'�B��svj�G���^x�lK��D���hȯ�*���>k
^}�$��� �!-�>���HV���S֎W8���W�y�����x�$��Y;+��$�r�H~c'�>
Vv� Ym�Lҭv�pxD��p�-k:�9bv�Ν�۴U"}��@n
)UUd�a�W-�+�>�f�d��\�W�0#R�!����*cF�xr��g�5b[�7e��o��a��q����]��7�1�V��:�UQshP�瞇,e�HǗvG�-}�d��T{t�K��0YF}�ue���5אx�t�^�|����j�KpW��+��Kipn�����0��,�:�h�k��c��с�����*B�_�R�C�r#m�JP4���*W��/�?+�4Jݙ�	�16Ax�:O�х���q�����������������=K��.C(����� �"bj���0Rs��� ;r������?�g�\ ��u�\�Z�I=7r珍I����}���2�>#�Uw�)�F�^p������Y�(�*e�?P�C.G|��I���;=w#ո_&�z9�X��ɒ�����j���}��>��=�&j.}��\e�:�!r&z���iA�!%��"��m1�v����Io�L�"�o�C���R^��=�';
�F��H^r}��$z*��R��%['_.=ͼ�d�"���h�gR�5�Ĉ�+ѐ\��A�BthL ��� ̊���XLv�N�B�,|/�o~[�;��(�eݜ��M��`$A#-n�hKe�[Z)`iJܤpM(��D 򝰊� {�_���,B�]�z�
t^m+�3E�y?�����5���[M�\{�,�v��܇�=댢� {�a��W�9U��� � <���w��h��J�vWDy���&���@N{	��
�JG��ޔ���/�֕ �2���\2���i�/��� �P-{'e�E�Y?L	�6뱔:�����;7^����5�L�v��>� ӳr����A �b�u?����.a�8�\��J�D��^R�~FsC��ђ0Jj��b����P��9]��X���)w]*�'wLH+=�'�݇���H0R�fJ�� �|¨¨������|�ȩd~�P��R%J�C����y��,ڤ�$�j(?#�iaA�w�o�wb�"��W�i(�;��a�C6�!�E�u��ܧ8'��Q�quj�3#g3uxL}�����m���a��_)��W@�Ek�cy�-F]�P��{��঎�t��F�;j�鞈D�%@ے��$OhjC^�$�]��jx�iqP>�4����Q�	,Q�sco�j�]��!�����HE�A;�&z��D��i*�
0QN�d�k�����c���H�����Wh�R`�������t�~��-�d�2����x��� 6����� HW�^�&g���0	�1�~�g�p� $��;Q��-�O��xP�Sk�J�u���3�����?�u�} ��1�؛��u+�u�guA�Dc�e�vΈy%l���������=�yU�͙ϑZ�}�h�G��kw2��v��!4A�K�J/7�F���l.ߐ�AΙc�����M�����E��+鵳i�v�z͇{�=�p�ld)�Д<�ӏ��2'֋&%�&�^8���cUo�ə�M<*��1��>��Y!��a�6r˲u��= ��؋0)B4�9Se�!�[�|��s���hl��Y9��{���:��	�h��c������t��YN�N�m��V�/$�8�z.��oS���e�QO ��Wci��~��nS~CDQ��ѵ˲T�I��!��L�yŕ����>:M����D�O��cU�36c��؟K��Qk����+OUI3%v$m�'�rE;{U�&�gֿ�h���W6G�":Ag'hv�r������F�?��_��j��>��Jn�Cr�`% ��跲5�n������Z��a������<w�I�z�ڪ%$�:��B��ʦ'�Qd�ٽ�1j��2W��$��{Nv��f|��DY��G���cDzP��?K����QF]=I�u�B�맀�Y�R�!
����?L��ɢ�<7�E$z5�c"��Rp��x�[qSI�B�jXF�,�w�j����A=
j����|Uf٬�b<��I�R}�K�	�?��$��3���T�*�����|>Ⱦ�J�����2�z!�����N3�к�i-+��a A�A.p�#����$�;�����*��W_��G�5s�ڈd=D>�mz�}��t!'3>���� ��7�re���vV���N��醄�2�=� ח%Yp�j��GLǗP�^����Дd���Z(�'1Nǎ�JZ)� �Q�A���`�M��E���]L	<���r?UeL#�6�<=}r?_YN 7W oT+s��tp�-z}�����֎�3R�T�=�b��b>�����t��w��jx�T�x+|F���\_�m'@�w{���:����m�rs�ٓW����eL�5b`�K�-���F9G5�¹���7M6����sCD$E�����⤏D�mpw02j5�}y�dO\��Q�=��ۨ���ϙ�	�c2�q�"�&�1%R���5~9�d�p3, �n�&~^A�p�|׋`�J|�����r�>��<[�R����t5�w7Qk���q��)��d]:�{@|��^;]̯I��$(wSv�]���2FtWr�u���0�j���a������z�n	�v}%<l��iK����)��N�5�G��Cp�v4����6���ܝ<�%��t��ww��g�e�L�ܫleш}�ޏ���u���۰�`��0my��EPx���`[v���W>��4�������Z�9\1������ρ�Jh�	�Û<ڛTm�]7��6?z�~�DKo*���E]�a����R���|��|R��M��]Uq��q7w�v�uv�!��S�sL�\7d@e�`CG�osg��v03�����������_Y��{�D���6sc�DB��/ۥ�؋de#+�X�Q#��Ӌ!y����ǟ��{A0"�1�V�ve�i��� s��r�i�U-*��u��6�Տ�(Z��ͧ�1g����#��2b�ssY]l�1s�Kv����;�C�}E<��y�����:@������P�����f�QP��?m�e#�[F"y��6�s&ܙ9;^w�=>��C�'F �.���~��b��
h=�����MT����F� ��ca�G�*�ʢ���\ߔX���Ī�����95�P�i� �l�#�����l�Ǖ[�F}8�4�pt���k*:`n"��0Pyy�����u��p<2�n�`�ѐ��
���?���y-�.�z0�J�6�U�%J�'+'�kñ��Π(����1-cSW�����G�B��j��a��:V]G�S�
ˮ�X�ȀO`o�S`aG���Om�Tf� �5*��j��Lb�����n�J�`�B?�QW*#����EkPMźwg�]�T�d�0m���-W�:�2� |���)�!�'?��n�\|�UNɛ���6`�b�ԝ���O��e�!&��U#TE5��cć/��H?α ��q^$e��hq�����������䐼�P�E�+u��.IZ^�<0��ݢ���=�Ю~uEl~X7j��#}�r�]��H�H��`�z���Ԡx*"c8�E8i8it��"!a)=o�`3�~S�����G�Z-�4�So��#���u� �1�y-v"����G廋��ز��ub���W9%=d��9oT�H��."=��
ϫ�߅��Hy��s����*��V��:��I�j�Ϡ%��q5@>�1�l7�	ۻ#�j�ܭΤ�nFa�(�_ɀ����%��
�i!�.+_90�x�(գ���E.Lt��-�a��d k�PQ�|���&��ӠR���GM{�[j_j��[���n��� �ͮ��E�E��'�Cl�Vk�eN��7>���8e}(ݘt;�\�x�K	ŕ��\M[���_r�P:�B��;=4��eA�yk7�F��LC.���mo�EW��8V�`D�g��
ήe5�9nM��~,]�1h��F&s-��'7)z�<���	�v���N��GQ�>����5x�Z�3��4`̪����8\��<��n�)�����ඤJ�q*�e����56�������l�$�J2i��SG����h%��p�
e�	�d��2�{4��)l�� 	x�Ej�Z#*��)���T�����}k<)-�-�W���Or��L�h���;��x+՜Lc�0���1Z\���!���)(�kc/%�E���c�pz�MŇ�?��Ŗ´Q�U�,<uC�DS���>p���h��]�����/��}k�/�7(�����c㍱C���0�9`~�e�@@E�C��#�~I�9�ƛ�t�t��W~0̩c�� �<�gGJxh�����h-���A[pW2g��ѡڬ�v�;��u�1�6ә뤕7ޥ.s3f.C§�rdr�6�������xL}#=�Gq�{ldA��F�w�_Y~�|��(��J�s�_�A�j��=��u���"o�~�����uq���T���"h�z�Yc�l]X����}X�lBd1���P��:/R��1�<R�������ު�a�Y�B���ik���ˋ�-Z���ݳ|6~��U����C#P4�b���;�@+-Q���9v�1��yN�Ӝ�� �
�B���,��ǚ�1��"Ӎd>�e ^���Ewl��`K�O �~�C'Q^��E���a�PuI1�EI���
�����j�/�D��)�1�(��);x�3��I�����N�ݦ��ۋ5�#�[D�Mb��g�9����L�.�I���xA������Ui�A����D��cڄ��i,VX�6%Ry~�ڏF���O�����_I�^㳂���?��] �-�HH]|���O��g����u⣣"������PJ&C�z�v���x����'^ho���y� Ӟ�I���5afE�H�s)����*� �f�FjZf�0�շN��A����oMc���(�P>)������58��$�`���KN�(w
U�'��H _��lř�8��)^���~��� ��,�]`���� 1ۤ\z�ŋ��%.�p{���&�R�ӄ�����r�0,`�����E��Y�W�]}ۥ���WBG'EW���u�5^]bRKl��Yr���Ww��	M�2)�l�9�O؈�����m�σ��a�r���é��6��.���y��e$,���{ޔ��]Wt_��ӒB@�>����7�4U�؝�)s��Y��[�C�\�%gm��#��0#P���[�(��ױ��g�^�x;���@`����<�h!�Ty5�P�v����!��� %�Ǯ��L˂Q���y�L��x
�K�Q���ND�_��P\��#�w10�M��4��Lc����R8��)�����zC��(j�aRh"�6(X��Rl�;�����x��`��g�|��)�<���?�]c���Ҕ T:b�?�$2��&��|�/
�,wtи	��i���7���[�����̙�6#<#�:�7�����&/�a$�MN���B�珫mQg��`���T��m������V
v����]��e�0-.E7��w]���QS�bP+ig�.ǼUA�M�33�Ka蓍w��	!�l��N�[Σ��Q�(pZ�e�v�RCn��Ҭ�X����ԨX���]���)�\��Я��v�k-�4�A/�c�2��,���roH�|�^S��{Kr�"��ǫ�KR-�A�hת친2�E%,��z���X�t¦�]��Ɵ1�Q�#ޡ�S�r
�9�B��j��ft��b_� �xv�g7r��u�GJ#�Q�Z;�T�%��ᢊm�n���-|�5E�d^a���-圸)����C
�������F6�J`.1^ã�s��F����B{p�I3K;�=���Qi.��(�Ce{�F������.�h����XG+2�wq�hYD��?�t����*8�`�y�nVOWW�E��'j�ώ�ojq�[,�i��ݲ�P\lyOd`���{얕ss�]H����Z9 e�p��7�0�Z���;j����P��=��;�~��9����
E=;c�����l.[�;�S�Ya`�1\�s��,�?q	\�ӨQ8�Ө��rs�pUi���s+碢�(E�������sZUe8�$��l9-vW�A�i�rG+��6�M�G:Kn]s�^��(��E����~;`�i5!i��%uD!�͛6�I w��*5rF�g�-E��6�K�?Sk�1_U�,w�=�>���rT�E,W��C&^�4��0�;��^7�#��T�do�7���t����,��\�L�p�Q-Ȉ���) =�Q9�S��\Iႜ�ʋ�����J���,.ʌ��3�,x{k�����Z��[K󈔵��Y:_/��:��d�L<3ϯ�����h2w')dp�l��SR���X�6N���Z-h�)����>i���D6���1�@���G�s�]m+Y,�uE��kz8�Cυ񷤀<d>��88���'�ϩ}�n $�r8x!ڗ��}5T3S�7]�e$-��$��[�����7De^�p��fy��TPE©d��I����j���M� eaN��v*���˼3�Z\v�q��ɞ�����@�Q�W������U�5�P�(����\�hgr&��Β��ԗd���x�>��Ċ\i��i�Uw^E��k ��i$1��,�՞r3�8�F^<�>���UݾX��A[�Hu���u�1�N�ST�u���/��[��n�����ت9ة:ws6+xr�qF��� ��η��%c�b�}�<l���H�����0ui7v1�b�,���_{�3X��&�k�Q6%[�Vo��w��ri1Q�!�K�a�Mֱ)B�9W��ֺau��Rp���6Q��hr�Q"�wV6�Y�o�k�@��g���ځ��cIj��]�|����o�����{Vn��="XA[�8�-#���֬\)B��b-[��䤁� {q����6�9D����8�	�x�q�Ǖ�M��ml��4>���)��[#��}חhPv.{ّ[#7e~g[۞��o*I~���x����q{M�@���k��9��rJc�k���X�K����+:J�$��7D��c����i�f����*~Q:���w�-���4<�c�(�y�:��㓺=P�s��R3�*˞���h�4ϲژO�x���%��,��;��J�Ӆ|����b!��E/}��cdzTkP��.�o��9��k��Py,�afq�=V��b�pMg��;?`��M�C1ا�r]qy���c���f?������%�����o��Q!f݇�pi���ҍ<[����G�^�Y�o<|�h,yreD�<k�<J<|�y��<��zh䜎��Jt	Y�e}�i��VO�Fd�S���B�$csMī�#�mE#�H;�V9��{���L4����	F�K�5���T��͊�cn-?ބ��Z��(j�j=pR\�����.VR���V�N�Jt@p��5PgAF�j����1B���z�^Kn޽G�H�>BQ���>uBE3�Lw3`o���O[��Oɭr�2����l{2/+V��b��@�ɗƐ�i<]e���i�ݫաC��i�MT]�#�DM��c5��y@Q^�n8
�����FmJ���8$?�H
��[*�g1cq�L�l8[G�7;g�g�R^���WE�����l��0��R06��u�����O[U�Z�vǝ�<GJ �/ +SZ��l%�t�/6u���<���q�\
�V�q;"&�Js��ZGRh�^Eh!�_6_��9g�����sv�Q�0��M�a�/��8��qȲ��* wu��&gM'���o�@��2�����K~q��`!��2u�O�D\B#uV!���<�������� �;��{���V����(� �wKW��E�ߣ��������w����u�28�l?ʵ���Ki��]C�i,�0#�=��M4����n�������|ҏ0Z?��Gb�7�%��ٶ��Ʌ5�X�u�t�Z�r&��X��ږ��9� RVŁ �0.
��z�a'��^9h�j�Bɷjs8A��)��g��i�t�O�Gꄎ�W ms�� �&�fM��R�w��`W��8�
��H�� �uC@���/���#4X����2fPH88��J4o)08RBYo�8AI���mcF���E3o�{��YOp��'|͟d6w9Ω5R�u���'ŉ�vj������U�P����-n�w-�L�"�l^Q��� M�KkdbPT�Q�l�p�&�&�(.�sR�~
���+ϟi['�ԥ3<]��J}��X�I�s�i�O`��!�u^)m�z�X	C���
��$�
�;��sGJbF@�u{�d�z�n����2(�Щ�ʵ.��A��nҋGmN��~l�X:�hJ1 �֯앯���������މם.�Y��1bߩ3r�H��_O���Wu�	�{�A��QG��O���;�e�\���O�d�ӭ�k�;�֎�=�?LfZ̺kB,���F�c�cOz�P�H�c9\�FTy=���*z'2^��:�9�/:8�S�V�'��*��&)Bp#�ãl�d�Yx
�e�`+A�(������'�5��/b�>�6���b9�^.�|�^8��mL�ܣ-���"ԋ3�dݭ�j�D08�:���3m-[~C�;�
i�j���
��������ۧ���Mi�G�	Y=�û��i0b[7�6�U��C6��Vd�Z�@x$$KRv-��c�j�K-��c����ِ��ec�Ӏ����ھ��с�[��=04�ʗ���	@&�hL�J��꾠ɳ;�9XL��L���h�U��'�0���|�����-���=�#�4i2ܒ�H`�Ц�G�rdg����B�uAȒ��T��>�^!���g��&��I
�X&��y�;!��yæ�
����V]I��2d~/��NY�T�uޠG`iGM���3�DZi����&�0��%��\ �( �U���cY�AL[�N(9[D���L��'U��ʌp�� -���D-�`N�IC[�M�&����u���G�~���|�ձ�õ����LG��Yڹ<�����RR����y�`�-sR����2���S�.�+9/�8N�B^'� �4���)!���o����m/k������)�����<ɖ�w�[�af}���	,:�ҙ_���դ�UPQ��a�� '�WH��wO��3I�2߸���q���j86HŦ
%��X�H�M�D�n~`/%��!'��b|/����y����_��?6T)x��5)�r��<�>�BW{h�^T22�1���Z;#��B��D��%�s�������ÍM?��d��rbt�$�FRR���p}�2�M�r�|Q���
\L�	E��i���qdt�����PS�2��V��5�
��#�i[���L;�q�����6�"�Βh�'�*F4�)yQ(9��,�xz�^�0�^*M����;��|�T�;�2�UoeU��O�L�OQ/�6���{],�P�!��Zm�X��
�Ys/gOSl?n�KGI~ޝ+B����[�'
�g� �_�X�:�vn}>��R����~�����vY�Su^N����;tM��?Yի2�ʀ���BV6��es ��]�k5m�:�!�H]����d` _jֹ��6q:�����P���D$�Q,/P<s���edǺl��J3�]'h`�-������-�.�V�v�*� >�^kF�;��`�H�d}.� �5P��/�%P�h^�0F"QGa��K�w54�u\L����Hj�/՘���m���HM����$Fn���%/��(9�%�������Ĉ\׍K�{��j�G߃����}b!�3�h�����
U��.��x���A���<�}�0�Q��rwXP�W� �����Ѳ��R�{K�_������klMk��~gvߴ�֯s�s���{)����Ȳ�c��Ns����'�PIj��Va�p��I�����Q��r�����]�C<t�k��:,�e�2S�L������\(ˮܙ�O��r���u�>�Ey�p�[��m,zJf�}b�'
ϻ���dG3�݂��}M�a�}Ǳ���r�*2zר�[y��V�#�0���=�
H���;�<���6����h�N�Ln���X���+~YWమ�NP�y?�o���Xb7���_$�VjD������hc��c�:��[62?�#�ġ��'Ff�>�i4�x]���xl��Ȱ�>�����)����֙��zɖPW��F��Y�W�Y^�4�'�G���ѥ/{�2�Ѣ9��&��W���-�𺮟����Xw%⺯+�]������"��$.�@��5�%��kzx����L�W$���ȷ=� �|�Hx�S�>�k���7��0�.�U^���e��)�����j^�!\��(ظ�o"e��+�L�va����Z��鍝��H�|��e�y/-�M����yv/��bq]��Xs�n��/	Cxj����g����Ҍ)�ObM��e�R��1{�t򬍉K����+	w�n��-�v�*��̰md�9��I���ގ o���8L�W�ZK������β�s�Տ�JD��i��~T�M��a�!���g�:�X§�"w�(G >�%4�{(TR�%���m�� �yrj��*���̘@$�ڠ�膱[4���o��9�f�`)y�Pu���z�eZ�A�:�>+
���$ջ��x�nz�Y�����L1�����xë3I"_��zL�i�'����k���Q���q��e^�-��y1�����k�������(|����IzM�k#+BR��c�m�[�/ ������R�zQ\oM55�=�۾��K�S�hy�����HbPH
��劣b�06�M���.�R��k#����>`jX��G��\aWN��T+��Đ$��?͝�������T�:��?]p��q�u�h�?B�Ͳ��KT �`�i�z]2W��b�O5a�9�M���:�_Y�P	e�r�C�d7F2"���U����l ��8Tlz��oN>AgLY'*΍lo�m�a�.k����.r$o�|�e��,QqQ,�a�;�h�U\�1�uo
i����P�R~�,��`����+���8����*��,��ML�?�6V^�'�3�����f.J���!&.���n.��Z���<�M��kV�a��G�bD�Q�zE(��k�,�U
���l�S�czŀ�����������:��tV�h�v��ʊ�=�,�B�ls4��u��6]�{���ΐ��-�S�FՆ��P?:�uej�:�9*X^q��Ǧ�y4��� ��O�.��vf)$��i3���g�k{0!c�݋�}�Dg]Aqڇ�L�h?�B!��m���d�lu��������FM�j�Pc�hNS>
t�W�2J)ג2%�k��--��ͱ�_c�ѕ%G��FK�0�s2珻��'�	�
�!�:�����{�*s;bN�  k�K�����ȫrLB(5�����Mͺ��E�Z�o�X����'��`��T!x�ux�Xee.6�p/��c�'�x�����)�$�H����hֹ��lE���T%���2Jܮ�h�����N���X>w�&30�b韯���ĽS��࿦��8��V���+�K���*��İٿ;�d!#僘o{�{��2<e�<U��{f��\F\ƨ�?��D�jO�a�)1�F�D_'�ΣV�������g:O���m�:�O���޷-$>g	�d+�VDR��)/��ħ����������Z٨zįܑ�aٚ��2hϰ�ZI����ÚF 
 A	w����� 4��z�Ut=A=4��\��,�`������b�!^�B��h��'���9�HJ�������< �����Q�PL�T�������E����� ��}ef�����Y.��:l�O'�Q8��q���S�d��L|PT�XQRu�0�C�ܢ)q���-V?���h����Q�%4�c�P���R�w*�'���ka�A��4K�h���3�����ҝ�s�4�@o
�F�1Y�E��C�A7���Li5;�4�&nK��ć�o�k�797vZP;J�x�ల-a��������&�eL�^J|�yVv���Û?M���8gN�Z�h%���b I�<�?����A�&�O7��;�K*B�T�?��G):�Y�d*�{��{SSP�5�Qm9�]�A-�� �-��,S7�b���V#YbɾNN9���=�ܩ���2}#�ޏ˸��Y>���<@�i=o��%�	k>X��"f]
�M�pty?Q�G)��#Wv�e�����\���g-YH��O>�+rլ���&&����n����m�:X��Z�Ŝ1��_O����f ֐�+��P웒h�9$/�����ؽ ��@R��j��[�8�O�QꈶC��_K�@�<bmy�{N���
����k7�u�ɂ�N�c1dH"Hb�D��U��=,�ё
�SҨl�ݞ_�ᣈ�+^�"��jM����=�'.���mè����!)�J2�[l�������������A�����F�`d��kP��l��b�YS���e���_V�6r7�k�r%��.�Ů�@k����@XE�QQ[8����
9��l�3��b]j|�a
����=Z�-�2V���W�����h�X�2��L�9;��?����e�Pb�
,"u�O�?Fe�7m�%
Cฝ�d*}� ;Jb�F�'+:��<�^
��K�ެ�������T���a}D�>�Q�b�](ܹ�?gB�w=�6I��ţ�n�:��F󊕲%�$�ds�K�a����Ai��豟���ۓ�CO���W���%t#��#^�շ\o�C�`%k'�Q�\	q�m�.�dmN�\�e�u�2Z�8�������F�?�o�[#U���r7�6b���r�_��O�#����^���Zm&l	�@z�7Wiu6���I6$�1��wp�&^DR��Jc�A�0����x.�`+"�9W����<2�������~�?R����dY2�KJ&1 �O���57zY�q(쳇d��ŐĴ�&�-Fk�|���]"5�&;�z��&�%��@�)�R�y�F��^k1�/B_<߅`��%/��<����f=Xɩ���-�6��b�")t��c�^��U����Y�������G�^V9����dٙ*:�r���g�>�Y/
�n�hZ�1�5��+���-ץP�1
�L_�2�|PI�R��+W�u�R�4�@ڭ�h�s�SLY�sH�r{I��2N·(����	n=��ӏ/�ʗo2�Ҭ%J�����G�I�~�"��&L��=*/ƿ��u&�|/0���&V4Ԣ�5�=��Ǩ�凩p�U�b��Z���'�Bt(IB �V�D��nn���D��^	�	00��-7�o��)d��h�"�r��j1�`�L���ШC3�B;W��~�'g�@]�ӫ�o�}d\��CGΰ���j��l5��RV
��#��� ����8���b�0��*~[0�?m�=G��`Ny|HF�x}z�� }v�Ve����Q�#�R�<�j�z��Z���E+!l�e�u����H�mH���F��R��׫���+�o�)�5����ƣj�\I5L ��?@2�����J���1{���%��� h�������iA�C}���s�v	�-���u���{!3ϗ+w�>;=+��<2EO2�؋�I�����+��OmՖ%CQ?��$]�|��B#s��d]7$����G�@��Y/��Ўm!�g��,�ޠuj6x�`�2.�� a���֛��͹�W� =1��I5!��D��z[���!y�r��^�l.��b���������aE���T��-{3�R�g��.�G��� %�~�5p�8	V���:� �I �x��7t�I���zV}&B�cA����*�"퍱��͢�X���]�p�F@a�<�0�z��"�W�E3��1E��L���i�)w<��@(�����`����U��3���L��o^���̅pՄ����������)��V�ɞu�$�9'_���X5�	�3r�H̆[�Y�{�d�jY�H�uDh���7�{�,����k
t�%2�e>0��N�֖
>�<����q/u.$OENJ�'�\�	��y�\&�[0��A��&h�l��Q�[(M��eUi Y�5��U�<�b*u��+�{���1o���ٱjf
՞#RwU�!#������\�`�M�3�"����:Wnr��Òy��F������Ep�ܟj?�� U���33�|D����8����̻e�G�� � $�czjU��:٦�K ��L�(�K�(�/�	�/�^�C|��
�H�d�j��y3�u:���p�C�O�B��V,�M���?�B�u���5�C���+>!�ĉArt���w�l+��֡��~Xp"��e���1��+�2]F8����F�[U�+������Xޝ�'�-�܂՗��
A��f
3�2q�+P���Vr��O%�01��%c�lZ>o���V���p�Î:F�!�^]4���&u�5���1�6��Hz�q����[Js7���i'I`T���������"�����,��`��<�����ǃ盬�����>��"��T}����ӱ������f�[�utrж�;�R������;���k�m.He1���d�p0ޜ��Cka)>����1�Ɠ�AGG�#yx|�=� �/o/#ʡ^(�ȱ����8rí���}�%�}��@�-��w��"t�P}�za�wc8O��U��"i�p����F�}ä�C�2O,
��SS(�W��M���?�H]����6�\�n�٥�-��in��qr�����}3k77��ź�	w����n���B|�t��'���,M�:�#ܩ�/V5�nuX%E~q��Q:��7~:�o���:���2�1*O��qeZR^�T�h��-��I�	��@'�>,���$z�}x��(y��b�0�*˨l0��
��}�{��<MA�W�X!�3_�[�h���x2`�rx���Q�!�o@�ˎ۝
�b�\	5$��\B��nm�����k��z�Y/Xe�����ER+/,��gc!_;\�SԵg�%�Ex��=v��؂�*���^%�xkR��nn	��gٝ��覅�v=�c�����f�m��#��@|:[����EI?#�\���vv�Q�ͼ�ޘ��芄P�Lqgݪ��yw�$���".�a��AEl�DM�XY�)fD�EK�v�)�\E���	X:�mKt���-��U�O�NYU�������_M�YU��ҫ.���ԩ�Ɛ�;�m��윐��ƈ'e��������b]�, &ܷM��?~h8�^4��)=��4d��xB�E�"�dE`sa��T�gu����q�"�T�eE��G�kG���A5T�L�����?h�)�I���9tL���'[�0�HȲ�鱡�ȓbr��᝹�����G��'���>b$��Pxo�-�$/�avmB��9k��s.�5�v��ދ�!� p�`5��EM����, ����g��L��_1t��_	¤<�@��	�	۳������������@�$�z_;���?~D���D��VO|:�9ǀb?����.�|���R~=�s I���m����ݵ�E�8]�Zߗ�N���+�~vp��QE�r�`��f��r��������V%@�Q�����o*��=VT?0|�%ɿ$�L9���� Hm�k����@��	Z*�,1��z���߇�Lg�6z�����i�0�h�e�\)P�P�U*|�U�Ć�*�J�)q��Z���ܸ��(�=G���!�cmU�'j�MRE]��Zek�����F�LC="��/)
,pl0W���b=�6���%1�w�d9՜G��ٴ�Y��A0��*�R}:�*
R�vRZ�)\�9�+ˍkTZ����}ĥ9�g���*�;SB)K�f�4k/�����aa��S�i����mܶY#���ֿ�[��r����O�e��G�jO�>�Mq:�m��.��o����>�I����P�\��ә�~�^U�]���v�\�P5ds���|_��:���Լ�&Z�����T��ȚhOd��v�VlK�[��I(�|��f$ ���m�齢�y�B)F�(�P���d�>�����D�/���㌏e������k��R�ȗ��(��io���� ��X��y �:ZJ/�� ߆��xl`X�Z�	�ځ��eB�q&�����$%V��_8O�����0):�k澥����b�H�ل�1h$�)��)�@7�A���(��Se7�3�Qя���N&I�c��2{�Av�4�|�w1�q!6[0{1/USM����LF!�����jC���~����f�/��Wn���k�h��ؗ)��'�����-�:��}��e~�l.��}U��>6
��N�,�XnJ��u6�1��g62?�,���2/�4f�Ȕ�����ђ+?��2ZL�l�g�TO�!S������)���{�o�����3��nE"�4	���܄xP�a��z}�@Y���������G�qQy ��R��ԲP�٣q���B��^�sa�m��6��l�oy�I"������(�Mܶ�&R�YT�[��Ù�J�iT#�����dl�k2�b�:n��E����e^5����5n��~�7��!HEYҢBI��ZIO5+ed�vf���,�'�l�3ӱ;\��D?��"5�Dh�O���2�ܳ��º��6�A�N�p�i2���m�?!��WJ�9��1��p��L�YG
DA
�e(N���C�޺�ʦ�ҙ*�oJ������g�+~���&���_:�̂�7H���B��g�QWO��o{��ӯ���)s�����I��C:g�G{>|x�D"_�Dl'r���*R��L�N�u�j!��~�fx�f�^AEZ�a
/�W���mw�Fn@݂ �H��8>l���`?�>f8f�	ț;���ŵ@�o�rw%S�#�-�fюn�?(@Ƞ��)3�pgW�P\!f���C���D(f�;��/��1$,b��������9��o��q�����V���ː#TِҼ썄d}����a7U����=��D�Ҳ �ȸ�_@���q��I�g���S��:�	K��5۔��r�I�k�@��+aL�#@.iϹ6�ٷ�-ʴ�&����E����RП>�q��,V�hfvn:�Te��\���r�L�q���qwy���3x�|z�z�+�Z� �Խ�' C�J;~LJ��!�u���V�B�ǻ崱"�����&�CQ7fa-4���V<����E����r]Yߖ˼{�k76ƫ�-�GY�.���R����*��A�z��l;/�o8 Z��W��?��v��I����0����Gӈ]3�M��7�m?���$��h�Y�3WZQM;��/�d��ۗ��F�D._LG�q7�
'M�'ʺ2����`nM9�I�df8���d�*D
�l�̀JM^,4��]��%���m�a�*4Eć�CI��X��8��C���V �m#\?��#��#l��Cv2��Y#�y��+���@��� �cU+��?ve�>r�|�E��g&�ͪ���·�D�롏2ؖ��M�?Qc2�r�p�)#�ί5W���O_^�k[�
t���^\��>WC��ԫ§�C�ݑ;�4�^�f=�1*�·{���0	���(�n��꾚{�_r�I�BzA����>�y�H�p_��R�K�a�D0�5���1C��� �/�^&m���U�y�����V+0[��ȏ��#���Ŕ�ݎmjZ��$�k��M	��� N�T��>p�T�|L�d�6�l;����,�6��I���׉A���������`��05�b�̔X>�r�܅�5�P�C�>$* v�`l��I�4X5�e����q�@_�"���Q�;>5��V�'!RU�H&�TY)��vl��b��3Hf2 �4-�������;D�9IΚ�l�z�!��D�ڄ1o�3�ܭqL����_,z�)��%}_!߲S�nUj�=�꿕KX�p4^&3VR�1T �Z�X������ZD�!��
m�d�䁩�z'�,�Ⱥ��^�z��p��]�n*�My��M  _����6ȢQiag�w�#F�0�[	U�$b���q��P�]o��ٰ$~�<wޒ6>�)��ʹ]�*�7��/]�����덧��Ш�����IY*q���ۺe-�|gDT0!@H$�q{X}�����3BB�W��&ʰ:�;7Z�H����M������{@\�x��0[��&qܩ1S��TFV�SKj+x�k7�}{"QV�,w�-��,<�s����[V��7ެf��t��CNmz�l_�����`ǳ��� ���R
h<���!5��p�30?�<1\y%���Y@Α"�NY���PX�H�e�ꐉa�!�^�3l��h)b�mw�sHѽ�\�SЯ���y��a'��&:�%�F$Ou�\�X�H$�`!5�'�ev�m�%!9m���D9\	�7��E�M��o��֨��DՋ�mLWa�ٌ�12�L�reA+�/9q/^GB���q	��[VJ�!�O@w}�o�&�D�wr,��m��CiE�n�����Y����\�I��� �
<�8������4xݾ�ZǓ�\ZژJ �^����9��Q����B2��e�|`:KJ�l/�[w�����T	��\Re��+���Ģ����N�8�(;X�p��>���+:_�2וh����S-�[c6(z�B��8�~%yl�7*pj�VA��f��ѩşʀ'�>pA���� �?^9�XZ�����Z���3#��v�F�v�8�)pN�l��So �@ ��fC4!����<-�L�I�9�)�ĉ?����X�K�J~�Cbf͇ļo��.��n(��L�]Я[!�h���حH�rlӛ~LWk�1����.��Z�S#�et�$�,�K�L�O;�-��KV��؀c� ���3[t~k 2uO����e�sH��9�JɁJ��������ֹEM���W�R�x��K��u4N4�-5�6�񆍝*mJֽěۧ�4��4-wt�q�ƅ<��V��4���'2�[��h��/�fb���*d�ٴ�;�~M~E�mb��61��<	��z�gE8�7W�x�)7����H��л�����d�~�l����:�h�,3�Q�oGN �ۊr�R%G7���^0�P3����r���c���\��*:�Ј��E����a���Pg�V\E����<�گ� .BaLo9��l�0�n�*X��y�R�)?����q,�73XW���Ɲ�[���q�f5p'py;��u���Gg�Ǹ �)čP�D*�h[p���%}*ż]���5���9��Q2���~��m�❉z{�;�A��ɜ��d��G�̓w�T�����	#�
 4��oUQi�?�=�%�X.��u��0MZdVE��@_����D8�=�T��\�l�Oa�6�E���:������,�%�Q�0C.�"�P�ԍ�!�T��_ʧr(��\؆�����EPL�`z�HAk3���I*���I�Q�#�x �	)�M-�7�0�9�}2�Ȩ�m£4��{�9� ��J�4��\��
]�W��
шc��Z�vS�Ef�� E��ĊtH����{g��ͅ�7�?��&;�.���,x��ge�E��,�����p�!�;!�`��O�ߛD�|�Z���Gfg������i�B��~��8��oU{�}M%�տI0�YN��X����)C�ld��|��=(��~�y�ĕ�q����ښ�SA���ZD�i��E4�1�� ��a0=ܾbyL���xފA*��=�	[$�:[&"��.qiՆ#X븆!�&�8�/H���XW~���{�)*��]w"zib�N���8��H2�Q
! �[\������m�A}�S.^�4��`&n#�,8��Iq�A����`��1uQ�����4{�PH~������F�.�2�z5[h�ل<-�<;Īw�U�$h,)�B�|Q"�i�/�:��t��5J���ǋ�iQǬ���_u_i)�oe�:JJ��9��p�4���%���<B�0�b�$sHz����1����<]��C�ʌ�I�`�A�	��([�����S��(���W� p�J�Lɚ��^���yԕcتk�.��.�`C`Z��>[�T���Y���D��ja��}f��� N�b$�)���p�-[�),|Ǵnz�7 #��N��V���p@�?G�l!���-2����n�l�f'(�<���8�lL���o77/�Z3��s��I`O�1meYC�'�XL!R���<W�3��Q�!c6�� %ձL�!i�tb#����-�k6v)�����]���C���p{�0��$�i �;��l������[a�5W�Z���m��c[#E�,�����~��������z�L���h�X�tLW�<C�"�5CG�� X��|��`g�ij���%_��̱¦�$�����F{`!�ڶ�َb"��Md[	"		t�>���r)�'z�����i��M���Xq������"����IG��r��_�Bo�`ae��Z��s��~�X� �_�_�?�._W����`�<�?|�@$�<|�Á��{�������(?�q�%�
�c������ֿ"��YJ�.�ZZMhx'��e�'��Tj�0�o&�9w�3ѳj�>S�χ%�;��"au��z5:06�{�?�u�08�O�'��N0v�O<8��������w|8��#R���:=(���k&���
����$�*��P��z�g�ZP���p��7�W��WK~^]%����a�-fA';g�	0��\�x��äskN�~��ݤ� ڛK]8����*�k�x6�����
��	Q3�ܮ`�Y3�X��o�͠�sh�A^��H��v��y[>��dԫ�(���Lg��@�\"�y�^L�Έ ��y1*)u�4�1�7b2�r*n^h��&���O�Ut{�#�f��c� �B֌���GsKg3n��4/�_�t3ys�7}�*�ځ	x�����6w�5E����c���Zo5WT5.�F��=�����&��7�Qa�r����LM��C ��dL#�Y7��G�k��ȟª-��?�~�w ��^Ţ�۞�ۉ���| }.��SC��ݿ%n;���_���@A�k�'^{��<l^�"�To忺\����:�e�)g�2y�~�АY"E!�Ǎ��?Y�g���z��)�&h��pۋ����|�0ua"�0 |��{-��M�.��R��|/E�u̝��I�s��}FJ�1J�q�`�[�s&&z����ku-=��������sb'���O�c�.w� ��/�Ȇ���������z%<���]�P��Mҷ�|��4,%sԷp�;�d�Ur�����D$��^"��;h3�P�����H�;��2������VØ,��A��0kī����a��B�X�P�~��\{�[t��`���+�6h_�k�jI�6J9�Ǐ37�y0��:@�-�(ග�E��m���C�e���a	,�P�>��Gگ�ԉ�s;�	rC�D�]�ِ�W�[�NM��<��Oc���B$���!i���� sԷ��M��J������q�R���(-=v9YG!;g���P�g2�#=�T�Q5�d{o�;��a[�-�0��^�͑tnM0���o����k�(SoD��  �<&(D`�LՎq���K�\
@��>A�P���0��?��[���'��שcY��ן)���� G$�s�U� G %A���&bk����$�N�ū��I��u���A�bI:|kM�`��dG��O�|_cAy�>���a+o����PqC��L��Ef4�>�z��!/Aw�����ױb(!mg�x%:�Y0������"��� 2FeM��_2�gꬥ����c�s�Vq�6h@OE���aT�	e5}�Z��(g��舌y����~�J������ )½>��	A�>_�Z���iY�:pz�#��Mh����q�Y�ކ>6)�`<L>�=1�UaE�E}��A�h'�^"Q��zx�O�g��	��P��-^{����^�<�H�g&��\�`fȍ����I4� Rzϲb8�Ʀ�&T�GY̻O����IX�(�I1H��E.'1U'&���k͂ߨXF��;��0��'��;YAz=��O��]{��-Rj@�dN�d�a�HU0�e8�O鯖�!O>�z�k���ENo�y	��g���h�c��2bh�c�DLu�KX�����h5C�P8�=��K��A������_H
��(76a�����ᅄ�WZٺRy$!��%ݼ���c�}�(����w�l������� �f�R�o>���n�bEA�Q>�}v��ÓZaTB��b��2Y
�_"�{6�����/��諵2��qW0c��I��cF��2�}�7NF8U��1���Q�����P.��m��gJT�mP1|��>�7(x���ޭ|��K*����N��^�տ��ͩq+x�A�=rdN��ӛ�"����\V���W�U8v*��I��ў~G��}VGnW2��;�s�C�ݕd{�@UO�Gklu!�~_d;��tuo�i9*d<)(�O�wg���>�������kf/�+�X����~�̏>�
wH�v �������;�q��f<���]LZbeA4�}[������3�6�������`�8�
���L�2����^��7 J|��!F5���0�'��f�r�p%�\ �.P��t�֔�\`�]�U~��Cg�x��g{Sȫ?wK�� �������y^'�^,S�g�M�m GKϫ`���W��2��y6�Cڡm�`����Jߞ�boH � ǡ���aN�^��ޔ)r����]8��+�/�#ҳ��w�G��LT�j��<��ǝ��z1��8��׵�I�s��1昻���d�	Im��N�K�9t�^�1��B}���CU&�x�����|�mѲ�O�����T��v�Q*�	ݡ������O��&��:����^"pe�t�S6����ױ:n#2{�3Y��]�ٲ�ߒ�~�u�:u����f�Hlfe�Qk)4ZG�/�T�BLI�B�o�'��@p	�h�$�8k���KT�Y�_f$�����qp��,[u�oJ�KDS#y����K1h�}��|�ZS��ƶV��.����[�-
1܅��h��3>��Z���v�Ձ�o�b���C輦m�/�ENN��[�~j�X}�+�Ҝ����ڽ��,���L1Lz��7o���`|kt�N��?:�hI��hϭ�`m���(��><W4�JFLf�/����/�U�d:	l�b=き�ݛ����B�L�+�M�}�w+I�7F$9�ԩ�a�ް2�g����M&������t��H6H���#�S	��C�T�̈ /�ȏ�&N>�
Cq�;�����>T��#��\a�М�V��S�c��N�Qut
�O\�/2���5&�v����B�[~&ۭc��d�2�J
�E��t�9�����jE��f^�/�
���kC.Pv[U�c��V���A���U��c9	����9n���x��H��rA{��9W�m��������B���|��V����Y���Ɉ�4L��
#H�qs�LU�GD[6՗*r��
̂w�Ri�r�.IM$����Wug���-*��>�Ʒ�HYbE%s�d�~��X>��SZ�#�c�澔�wO�Tc��!�:C�E�k�1<��i�u�"Xi���Lb�Χ��/����[&\tXu� pѽt<�+�q�A�:u�6�ar�7U���'�^����3��+�k	h(Z��[�Sf��o	�`��4LS����z��=��Z�Pde�Tu�IO����_Ł0Re�%����7�Wz�$������s��zv ��&�@������,�L�����TM�Y-���}�$�~0����; (�u����������F��Q��]�諒��Z����7�r!Y���1;*�To|jkNÅo\#s��������ov �.���-"cA%s�7��{�\�x4�0�b��*�0�@VOK]~��uU����/����ݢ0� &�a��T�"Pe���,ҩp��8���LB�#��?N,�Y6aB�Sr�-�@�gF��˟���A�i�&�hA^�4�͹��~y�1��y����n�)yIh�SHhC%�������}cΆ;$Tk�~�҃�-���_�l'���OK��"j>I��kt�����9���(��^��&7��;x�d/:SpYI���h1�+3F���?����5�!K;$?���4��n���Bv���c��;���{l0��+�[�<��w��&w�K.���*�
�r��\GR�T/�Ys����g��o�!�_�4�/h�>����"y1��x�¨�2��ճ����
o\ / rzC�gJ��@�W���W���KgJ�vqQ�0��_�@�
��kQ����+�Q9��'�M}��� ���5����1穝?��뜂*������l15&%�,�(� ��۰>L���P�C��WA�k����A��b�l�hI�q�a�y7:J|�Ku��F��Jr�8>$#~9Ցx҆�-#V;0}�k���#�{*�w���}u�]�����(�Ć����ȭ=��������`���Nқ��z��g�B����m�DU�n����m7�!f�H�	��2"c�F�N�s�H��s�����z�gew�=G���x�����}��^��@���	Q�=����� �Ջ����:��BpT�$�� ���4|$:�J׽�aU�rT�]+l��N�;]���Vd~���p�틵q���[���T��/�|$�KxY����߆�r���=��z%�lg��<	�%�x77�[��t_
������T�jg�ic�i��줕L���@��3�$CM̤�izqr8R�tD�Ł���,g�"Y�|!p �gu�����j2P����uxI����D/��\�M�w���
4�Dנ���
+���1-x���s	,`]�c
AS)�V�C�'����g�:��G|�	�0�^���Z�T��R��L^0�w2���!�5�Uy�㱓`0�ЖpՋ�,t�h�oc�4����:7'�e(��@�G�X�iu��#Ί�z�%����.�	�K��b�0
�6�7�)R��F"��R�Y�Im����9��M��gCL���À�-�����QԚ��Z��^�S�>���GJkwO$z��tn�� h]jڌ� h{�oj�Ɛ���OW�La��og�~%��Y����VgI�ۃױ��L�i��?ƣ ������?~��u5<�&;6�y]��E5W��7ϖ�bֿ�����HO`�ɚ�aۍ��8~,8|�Nߴ�ʽx(Wqn�P�N�@'�����������!6W��; ���#����� �e�a)'7�W5�p�Y#�EU�E�S���{\��Kn��ӌ��R���a�5G��#�.#5矪��c]C���k�n2{R�}����"f�
�ncO��@�b�}��	`��V"rpo���{�����NC�1����K��s���"�<�Q�Q�(1�J\c�,���Q�*�s��
����'j��o��T��/�~K�Q	6���I�)qZ�ŅfYZ:�w��U���ٝ�*��s,���
�`�pɲ^ݪ�t��yܲW�LW�^����	�i4lVnV��D!_S��¬�����E%�(��_�q�+8O�T��.@��A��꿜�C��q�U�u��r[}���L o�ۄ�ͱ��������J�v��@~-z C���_�<�w)�j�'��8$���Όnu\R�@ J� C��$;_���rL�"Z��+��_�C�����`���u�$y�W}�哤�%���O�\�=L���`.�a��C/\�;��!��"ǁ J-1E� *�?,H�\�˲�[��2�V�R���* '%�[�Υ�d�8�]��kVC�z�
̢8CS�=V^�ċ�3E1��}>7��a�4�r�
�ۦ׌�^�/��o�%�^�P�]���/)��z%�#dM�K��ٗ*���^���
�0�VR�V1�4K��J�a��",�m��w�	�3�@'�h~��Rv�_��[�Y�ذv3���'�
��Q���ް0�9)��H���I�(8pL)[�s˚������t�W�DG�ݰ�p�Df����LK��*Me�Q
z1�k�ф-�N�_��2�Ѣ�'GQ�����	�������#]��,��)(E�'qկ��K����O66�I�����y����R���7O,ķu��r_cUz3�A>�Xs��I���s�\R".V�mW���ϵ�BJ����>�{X��E2!���z�8z{���JZ��jF���͚�V6* @��O.w�"��$���,Ӂ���v���<�ubw�T��0����V����A�ːLC7�N�	r��.S�x�:�0bɗP�{��w��'���"p�;�y�=&9��*�c�ިQ���^�Z���X��AM�@�UWҰRv� �|�M}��&�I=�"�t��셬;��=�ȝ�5�oo2�˶*a"��@r����l�9���rSq]����5н��"�L�\9�N��ӵ��F��o�q\�I�4L��M'Qڬ37���D�3!)��O3Jk�lQ�r��F�����W+�P�u>�B�E4�U�[It��ྩO+������ٯ�%R	�m�S]�?��)f�Q��ԗ�A% w�m���r*��Y`֤%���jn�t1?U���[��R��t��cII20:��|m�u��M��]�f�4�k ��>��ęf㵀�(&+���z^힅�Ÿ���婱���@���oa��Kv�*���Ig�4^���*�QtG"����h��U>9��Y�O�n��6�����D@T�?���^��,~�G=$Ǎ����m\ N���3����9�^�&$�x�6
�����5B��?"�5��q���� 	�����p�;IԐ��He :����}��,:����Y#��������@ɉ�Q��+�0��&�I�N\�%��{+bݔ���sr��wl 9:Ԏi��dƤ�?SZ휚�eJ	~��]�&&�"��� J�BR���r?P��Sȑ/�}p��sG��7+4�׮���Y��$.e��#�)�!�����i��QN�:�80i�-J%�(�P�{����`���K)~�ň��^ ?��-٭4���	FZI"��Z3}ڏ&'��N�ϑ�=�1����I��'8�fU�%'�-�UjGya�a���]'��J�+@r�0� ����E�~7�#B
�s�f�4�ׂ?R�t5���OZ������U���ŕ޶ f�ޗ�a�E��b�c=_My���v])�ԣ��yi��O�!� P���3ű��`�2q�kY�ړ�P9��m��Ȩ!)��G���S�k� �^�d�B�0�D_��|�WSFu�T��4��`4/��j��Y�eT�&�(Ʈ,�o��G���L���13�3� o'D�2�[����1~�.����\��@�]a��BL{o��^��M�(��L��?J��5c��{�>�����B!f"���ʩ5ݛ�]���!�0�)�T5-�qs��>�� �5`2��G&[��w0X���FFbl$�u���r��d;MC���ʾ�Iyg�U	o�x��U���UP�^�L�K�JH�}֧-LK�љɇvw��ۀq����'�1����)y�!*}'P����n�b�w������s_c��?��ʘ��]Brb�_�wf�,?	�� ����'a�=e� ��u�PE`���s�N�:vln�c`���J�mR◴��>b�R��d@�]Ƥ�:vD�}�o�E���e2<�Cϣ.}Q��R�'O��n-��-�C� #���o�y{[�ƫ綽�O��(�,�������Z?68���C�'+���i���֦e2��T���"�Û���՟=�<>V���������C;7��i)a�M�C�.����FC��E"i�������W�-H|�"߸.R�}���O��iM^yB,[�<�[Z����U�I)Zg�A|���Z7�$08R�m_^Đ ��$�}9��X��P�NhR�ؐg��m�0�8����.F�F�e�I�~*�:C.��%P��)���Rzj7��<|��8��#�#uSU꾩�^���"��%r/�%�h��%���'�,�7���<K�&��G�]F=���S>4��/����JrN-g,�'�_dXڪ�(^�菧����6fΕ����/%.3���^;c����<q�1|y���3��4����b�҅�Q'�N�,���5Џ� �fR~�BRж
�s;-Nn h��4�Ȃy���}��K���T��SۗW��8"�v�D��A��TcWn��=�(;��� �������v��oA���pa�>�墳?�Q����}2=���v���^��oi�e���7�j�?O,�N,dq����tl(L�g�3�i�8����k0vn`M�/�oXD`�neR>F�^yR�{4�=�ve����-B ¿��ПK�����ĭ���D�)נKO�V�/�j\n��,����1��l�kcR�N�*�}�*|��k�������P�ࠒ�K�|�<n6VÊ��m�i��׍�I�`�\J�ꈄ&}@s�`%2Q�i�^8����}dH��w�mA��jë@����������p�M�4(�@ƜcNv6�{lQeP"�yc�z6b/(峆��S����y(�ނv"���_+�
�{B��H�ax���5��ԅ=N� s8�J+�߽� 	|#�/&���i�.�.�fs�װ��҂N�w,0)��qU$%CҦi�G
H��E&sNO�:k$�����宓��Z�f0lM,�\ @��{�-K�Nէ����M.(�� �iDŸ���AO1����o�"����9)}+��zP�v�L�4�;������⚦	���,�:��C%��pd���pA[M�"���Á�S�� �e�O8�Bܩ��{��j�F�!� k��Fc$��e˅TZ�����醀5���Lu��πj9䂡�5ԜA �.4�@�|�lT��پi�mi����A#���8���'WB�9��C��56`,z��,Ԇ�?�w�l">}��4����)Ic�(�u���v�5=s�
��L�%�]Ŧ6����*{#�LX�s(�aQ�[�Xl��Cb�s\���Gq�sU][M�/�t�cX�;nZ����o	J�~�ng��g��CC'�˶�ߣb����^z!�̱��ZL}Ԁ�y u _n��\F�֫-o�J׫���
���N�'�.�&\R� ���jή���Z�qZHh3/�p�vֲ�T��*���5��F@�D4��&�KK�kq1??1h�^o���H�VV��]N�O8H^[ﳴёb�at$�bb�o�Py.�%�m<Ӊ�"�C��]Sc����8Gh��.�x�x>��_���u�(p0ppz�%rB�eݙ���� ��u��0�q��B��٘�UX0��/m.ٹ�H�<;��J�=�X�����DV'19�Vب��sm��*�4R�a(S�����
�(�jȈ�}�����k�&��E"�S���9�/F��~B	�j���ݑ����H; 6�iW��v����)Zi�u�#�ZH[����a�ׂv�#]�@����{��|�l�����ԍ�&W �n�.��0��~�z��wv+��
oB~}��ӽ�?ύyHp�x x�~h�vS���?&)�2��Gʴ��C{?U����2Gr]��e�u&D� �\ ̳[�	�:}�"�Ȗ��9<��~�B�߲V���Jv!�����䋞�Т�[�raz^���w�XH�%E��v��N	,��V�q��6Ћ��ͣ�Į�Z�)��r�H���H ���Iα_�o��6��)�pp��o�OzN�K
6p�?-u|��@���c��'�tB��~���]*��K���y�f�C��F^�v���ji1���bm�qN����S8��2g"�g�ۄ�5��i��h�Ɲ%��1�1�Glc�T�_I?�]��dl9���~f�v�]q����r*~J�ЈT� ȼ���{+oſ�q�<ֱ��è�b�� ��EA�l|�_���Ш׆�y�.�����z�/�R~KK���YF9���� ����5�6럟��$�/�;����}b����@�T��?b� Eᡤ"E�t���k��O�1kLj��qeW� ȎQ
5�$/j��D�O9�w�Vt���֑��@0I�����-�]�7�c�F�ĂK��y��`{)? ��:s��Q�767:E ��W��a
��ٞ��IQ�ߞ��C�6P|�=�bQ�w�w�Jl�U6�QN3*����,Ӕo�@�;� �>�����د��aӡ"�qe�6�E�\�%��'��[��4cӁsJ�Ӆ~�I�F!����B{�j�b.����M�����~20� r߰��.�g�g^6�����[� 2=u_��2�e��ʕ�d�.Bāh�zO��t��Zsc����L%�Ad!�Ӯ�&�*��`ϻ["��{�p��d�%0,��`����Z�ꑌ�����_�l�&eg�;�h�z�t%&�[�O�6��]۫�z�v���Elr�],2�rІ��bn�d�m%.���EB����b��e�LH؀t�ҝ[X��!��/V��'�?/|��x�J�s��Y��[l��ȐA���;@�����G��.������c��~�����h��z���f� !�0.���57n�[b�z��SF��$�Io-k�G���S�\h���"�i������P��a�J����P̴�Z��^/D�5=5��{s�)8�6M�R(��s��`��8���y��)zy�BM��
�W�5��������h��چ2V8M�;�^R�_vw�t�0G�8֌�L���Q��D렂醋b�M{���L7���g��G���������t��Œ-J�&���(��?�CP�:��������o�5�'P_$.���:+��L�
+�l)������w1�E�m�c��J�k�(ވ���k��R(�l7�9�f]vR��Fm:6�\+���ݖ��\)��M���Na�W�m����f�]��f�W�$ue\8������Et�14+���æРEڨ�E]d/�X�&�O��]S����-�9��1��n��đ��n8��V��?d�%<�������ƯM�4��:F	���S
�7YK�\���ۮ�Kgga�2�Y` -ΑI�$H�b��14��jM��d��2ϒ]W@��ns��{\��l���JCO	*U������%� V%�Z�lSAG���fߌ�L��G�4�z��q��?)`&�-��+��e�W�A(���j��D�)�-/M}	V�:>�jH�L�Z�aH����I��n�rkfR�#P������Kד�ˉ����1�A(I�ArRoXWO%`� ��z�ZE1��\x����������z�LkQ)��V����rүM���3��E���|�8��*��w�����K�/��(�y��-1�^�Ãf
�dƫ)�0�Ϝ��Ue��k��Z���*n�Rs 	�� eȢڱ��h���&T�N�:��|@�/�z�60lV���T1�p_t�#������P�Q�Àh]T�v�F��ս��$�@J0JU�.��Z��P����p�u���䓫^�f�"{I�G��z�!S�HAnۛ�C�xPc78B�۴����&d]vw���Q�U�MFC�r�tQ���}a-L�j%�p&���jт���[@'ד���db=�R�����f��zH�o�����)�-Pw+t,�hA���%�2S+:*��{�l4?�l��eϝR��qTd\Y���8T�����ݠ�|75���Rw!�x�e�dy��o/����p��$�����?�(����2�J��ɐX��T�z�o�5��r��	�N�8[�i���J�AV��wl�Gk�NEG�7��� �e��Nx1U�����N��/DjS7�A��u��(�F��� ;�^HdْGw�l�2H���]��9Y�
���4�@߮�J�"�f����o*��@=9�f`�l���a��0nV���~UK�(�ֺhQ��i�G�*U� ?����W�q-��L� ^��z�2��!y��	�Bk�x���:ڲz�I��'\��To� >��~��4�� D(�>5��s��9��	���� 1��3EA���*�D�u�-�����L��ji��~8��Fo�̶3���Xذ\��ʎ3`e ���#��z1��~+�6��4�q�w��A3�g�sr��x94��Uop}�.��ؕA=�f�[�`�Ҕ�/������Һ��Q�=���]�p/�v�.9.̛�xa�т��b(/`"��>9h�n��N�E#:�C�9����Ų��^V�rh66AU���q=&�n�=�7���� ��B��"t#"G{x4��Jf%d��Hx!��Fِ� ���9��p�$�T>����8L%5"���C:�g��aY��w�A:�Ŏ�Y$[�8����^0t�eEB���B�6+��p= �_�OI��~��	ݡ���� H��YjK�MK�b(��#��Q�P�S��I9p�	8*�}	�-��q���N)��U�{����k~�B~8�#vYJC��Ѿ�����'���� ��'7�3.�����\�2c�)�|��f	�q�Z�&�X���k�X��3���1��԰�6�#$���=jI� �L����sU'�mԝ�D������6R�`��Bt�z��/���Y�󬨨�r2���K5�5�x�&�x�To�CE��6��m���}S��'k�����rg(,�y�\"��w?SE��Z�
c���>9,G$r}��ُ���Z�ŁQ�u�&"�|!���L���;�dӈX��vC���e{�%ǉO�9�?j�������ȱ���J��j�w�G �#)�F+.P��D�Ʈ����?�-��-g��1�3D;���L�uh�|,��e0Gw ����~����9��������������2�#2j��161w��Zz�M0ೄ��Y���@���^C� ��"p��7���?����:�~"s՞J��#�)��_�5{?"U�x��ɞ�8:��� ��W%^e.v0������U�r~����uǀL̎ʲ��9�z�(�G��"X$I��y�vd�m���`R[��QX.X!�mc�!�!��y�� �_�d�H�\I�
��@�T&��3��̛��/�g�=a��>鸩lkW��^<���\C`[��O@�k�16u��ܴ�P��[�8�|��r���Ϩp����J��]s�Ŀv]�`���*s�&8�J0V���MD���3܏b�YR�h������a��[S�JoS�60��Q!k�/QMm*A�#R��:�gAW�d��j�&;����ާœ�>"�$�|���i�h�oHš�p*��<�n5%�Ґq�\$9'$Е#�`���:>�'8��QD��UER���w*D���0�F��$�Y��-������faQ�'mR�ז�J����Ol�,U��R <'�� �K����OR�$G�HCG�҉id�Jhf� ��9�f5��y|W��p8��݌��5_U-U.��{�fA��|	`U��闑�Q#G��q�2�L����r�|&�MƳO}{�5�ʉ��^M�oWQ�./ �Q6�+N]�����i`���D�6�K&��s��Z'���e\��?s_�*�CЮ����?Q��Сzc��K���U�\ NB�E�F�E!�vS��[�<�.v�-�����ތ�*���K��װ!������dD#h�R{>��WS�pYY��L,u�<��(�XѢҒ�T�f%/�֛G���ٹ(�K2ˑ�>�m��ǫ,�*��;�pW;{?H�nR E(�R�Wh��� 8�pQ���}�V�� "�jn^JC�t��ƅ��kjwfv����i8"�ي�o�WLɿ�a��y�崁ͳ��m���	�=ƕR������F��M����-�����)5�RquY�yA�C3�έ >2?g��z[��^ƶ��豣�bĈ�)h�6	B�~x�!A9z��Z�B���O�S���j�k�?�����7^%c�Ԙ�	dEN_ߩ�5�Fp'�t���%��Q�Q ;�ev�ue��0ϔ#&����9��:�ɐ�P�r:_��@���ȯ�S���G2|q�:���ƳS/Q��o�&R�C��|�fN&�*���CRn���ĥ�.[�Q�'ei/�mN�)��o�nm�4�}���FM-���S�Qo�6^�b*�)N��>�c����S6:�A#ʝ^��j�U�.�%т�>4{�6i�씍3�b����7f�<T(ĨD϶�#�B�=��a����c�JTc�Q�h��:&j�H�75�C��Nffm.
��wp;��饋�ǘk�R����{� �<B$TSPb�G�v[��,�g�C�N�,������34Z������u$b��\ݔ0�3|D3{�JD}��x�
)��r� $�C���B�w�c��I[C�7���UFR���:��>$�aF_�Ȥ��qzݡ��tU#�Q��N��?�N�.e�S�x��Bosiu3H��e�����Z����է�C/�H�	R�q��Zo�����1���)295�u���)��3�m��W��ӿ�>�$���m~��[�h�q�FU����(^���a«��FA1ߛ-	�����6�{����FE|�>_i�RV����y1L<m�z���f@���0{ȧ���"qR�1'���t�3�+aF:Bf�j6%���:�]����ЙB�J���LB�Cy��d�*6E��ޕ���'w_:atO��a/�����J��u�X���{̒ʑ���삪����tO,��Z�(����Vy��I�6��G�K"X�F#���#8�^�m���*Ic@�5�4E����{�4U��\ �y��)���" �E�njz@��U�MF�

��Q�`���.��CA9�N�7L�lՕk�5"������s����tԔ"�8_���+υLV-���rwG��%�M�{,��.�������:�w����sV	U\:��6����- ���3��x��˼|�X��W���g�����"d��R��^�ZK/x�@�T@���.�H�i#�Fu���f"�.�����˝Y��f�B��i�ۃ����~���];�y_�(d�O��f�$��!>�"mf�$/�@���@�J&�W�d7�Se�Ӯp;=��p�&�2�VX�����ї�Lfb���Yf��� �`$�
�S�j��IunQ��:�DXQ�}Q�s^������x��� ��O�	#�Lub,�<Bx-�*��:#��[L5F%�%�6�AV�����j3��xR��S�eQ��*x�
�s����>o���ŷ� ��`�	Đ�XL��k���-�r^��/��	E+�8~&��p��3S��|���u�8�z��li^c�3�yQ�����e���ȯ������r�4��y-+~K���YW����m�B��1̽,�e�?>�D�`�侐����c�Dp&: Q!�MT�������%���օ�HBA�V p*w��ND�>J�k�&^��u��Xr���z�3i����� ��}���Ui޷O(엖'1�u��j�~쵢^8=��G$/B�W@Ĥi��+��;���<I�6�b'[���ՙꈅ$���E{:n�
�vZXp�j%��{�0Yt7K TqOq	�^&lxo��UU5f?������|w�r��4��^���HQ71CO;=�W�0��9�w�U�ƫ�"L��Q�P˲�p��w@�d�n�cȹߓt�h�����t�{�%��f-t�w�� .��
G�>3u�/�v�>�ΠV���o�8����V�$AuC�N���R�Y�	;��P9������j�����уt\u���}���[�9B��4��*1��25%5DC���7��	���S�Ԡ9��ß1�L� ��KB_GW(U77E�0��GM�u��,��}���\ \d.W����6�"�@]v�5)�J�=��?Z�}L �jC��zu`�J� f���2����zذ �k)���)��y�g5�e���t�RW�� '��{��9��_*���8]��Z��ja�.���޸mf�����6�CK{� ���CV������t��u�������|��䡫���F\�cm�
ԱM7����:沭mq��F�`�����f55�K��W�����ɏ�W)����7S�SP�7hs�}WT�3L�����|�M��1Oq#�	^G�Z;���Th�*��/9G�>9���Ƌg-��t�j����8T^�d(<��K�<��.��k'z�c���)6T�N���f�����0$lO{\Lm�������D[�k!ۑ|rJ�(����z�f��OI��h���j3N�"�ҺM�<cM��6�^�.�|b�1� c��dw�G��"2.V�v�3/��;��3Ӥ��;��%f����)P�?�c�U |NV����VL3��T�*Df�U��Bzװ��uvד"x�`~S�5�Ŕ��A�MK���1�(&���P���#N����);>c���d���r_�:ޭ��0b�{�p+���&�9��v+���/r����;0�ǎf����bW�d+���)�ٚj��w�OHg�����1!�Q5]ry+�'� i{
�ey�]][,w�5vѬ��� .)Xizs�t7�QB1��+�^�H��M����)�g:�4aT�[��ȅVWZ��m�Q5'ͅq�_����5�)-Q~U̥���|UY��c4�x��'���aL��b!�N���ew�'�>5e�����4'T �B��A1�F�ub��vo�svA������q��`���Bu�����_Ѣ��I!�w�S@L����� ��4
���_x�y7{yZy!�4��^ol��7��/����PV���_���؉���Ut�
X���6�)�w�q�;9yzLBU��ڟ(x���d*&��J��SK�#*�\��i�����������&^��`�9,�	��8�s!��(r�yaQO���l��~�QA��T=��|�+R<�\R4Ry:;��1[���l�n��p�YG�x�xs�=U�~`�����l�*|�@��)��̳jH�=F�_ ������jm5�Ӱ2�ئ�t���N�1�y��०9\A�& ���'e�9��M5U��g*'H�?���ʝ�LDc'�a���y�ⵙ1�?�%��쉳�{����0�5�?�.�a4ɲ�?56������a��(6z�ה�*�ӻ�|��Y^�kF��Uᕳ4+p��u�*:zPSH�QՐPb�����绦6����",�Mݠ�\��
��t�؇ꮫ�"zXg6�r���ڋ{����u�W�@�<�Az9eI��(y&8C�ȴ��c�2�4�_;�n�d��y.1y��"�^8`�h�hHq���IC���J�>���<���]�W%U�5�� #�!�'����7`��xOo8�n����2~b��C���?��gl@b��2*:�D�9g<�kN�o R"P���?U�=��ж<�����xsp5L�t�e�>�=9�>?��>o��_:�j�q��aF��齆
���%9��h��{+ ���M���X��9���;$�����v���V�D��2a`��	�zMl+������kʍ�!���G]�R�:��Ȏ�UB�ő-�Y��=Sarm�>�0��)�B�Hy�h(;��PV�]����m�R#uMaf����8|�+�V�#"J�@g�f��J��w?v��Ue��v��|Hb%���d����Ӂ�d�q�OV��T�/�\�D�:M�$�Q�ޘ��8�[x�*M��pB��c���+Q�T��ݸ/m~<�я�<���C��t�'!0�v�w�oԊ6��1�C<Î�V�$uS�9�7#x���G@����e���u�a]jZ5^���n�_�ZE�����
	/~3h�Zرbf�n7�>��`��X���7���4h*����#2���5��](���H��$�����z�����m�xR�}-.K���f�Rn��4E
��@o�\j��@���0��+�!����И������zR�d�g��XS�+P���b�m-�ܢ8�A�O��{�h�9/��g2d ��'	�F�1/%$`�P�I<'��
�k�⑊*��\�;'�������O��L=$m{��%8�j�����!+��Ca���$�ec������ a~�Or�@8漵��������&�#䟋��V�aB"����
�돟���嫛W��`��5HPL2+�:Tڴrl�~��qs��`����"��HG&��i��sAb6�/YKL_�`�Z���Tx�fOD[3�=��,�P��T"����M�w�u���m��?��)[�ӦF�/��ZZ�W��".*��V0t�ԝZ�K����!�[�g�-Wښ�*���-R�\�r66�&��l�}�-`�
��p9k�Є!��\�T^�9�Ѓ۠E��\'�s۞A�E�I@�6P���oC�a>��qT0��g��_}�zu"Ans	\*'ۄ�{�&���@����F�cMܼ{x�ه9�*���B��0��Z˵��s�6����/�65<r�<=`D��)7�6�S���}"�{�rMo��ry���^v��ʌ�pC�)��h����/'Q���&��W�<���f?�)_8�Q��a�.���1�D$����aT�����h�;����ҧ{�/�)���V�\�?
#͍�_q�L%1�����F]��_��J���>V��k狕�n�U�V������\Xސh�����xA�gnJ[ς0�A���u�W���8���tf�~?���qb{���D���V+^�����7�@��ۯ������q�����Q�B]������f�0Uh~��[\D�/�G�'wy��J�h�9�]!9��ۚ�+��E�\�-oa���;h�Ug��E&R��0ny�<�"��\�V�#��c����B��X�tG��q�7ث�GBL�H�<Ch���"����Nm��)בw[��T��17�9�٦c2���x
6��r�r��Ay�n[�g)Usf>7��L�~�fbH{kV��͏.����M�秮P�B� B�muryv� ��b"u	�v��~�����zJ�G���2�i\=�K_VӉ�Swwo\�/���hf�nYaw�LDK@����j<��MM��.����'vv1c<S�'a��H���'1y�Y>�4�c��atw�{�i�@է��5�ᕔ��ZߺH 5RDq���DT�^���5܈*��"���jJ�@B�h�D��"޽��oxPj��}��r�za��P(cr�Xn.%!Z�Q��;BI��1)�%M��!q����K��P��!�y ����������.�r.�Թ�K�n}���� �.�����4�K �����e��s �'m}ȊYb_ω[�P0"����`�G2���i�����-�@��RΗrՎ��\8P�k�"��K�b�.�7�E���Gn�u�u���3��F�hɽ(i�ƍ�+d1�8�}����	{��B-����G����눙��!Ww"͢�r�ꆖi�|��,���A�����n�	)�F���qxTBm���s��������b��V���_�ɜ�Y8��1�Ԏ\���t�>�԰$�j�d%���{���X���w�8���R26��kYpx�O��(Y�����w���&_�oOT�_ȭO��NQ���7�� oѭ*��*��ߦ�!ݯA[	Sl�����u:�ʗ"����eAJ��;�4qM�Bɭ�%c�"Q���C]-a�9X �V}�s/�7����at�t�)�s���¢�Zqnh�Tզ_K�1���uc�븾����Y��9�o$��M2NKkK�L��1x_�R��
��*�#o}�×�Ҡ���s�o���0_�3�TUW!�����`,b�y��u6aa�a�9��0�;��˝�D$����+z��;�YQ�|3�y�N3a�3x�D�O�G��E��+�ձ���ó!b�{Zz/q��򓧳��`�&�|��L�G�A�2^�h]�l�+C�hRk���lOX��QDCX�z�&�CPF�-�$PIIX���Q �B�CA*����C`pe4}�j�S�	%��gÔ�uz�;�p܎O�ޅn�Y��.ݥ�)6���ϷAU�ˡ�Xz�ķǡǺ񪔡J�ȁ�.y!�nSP#��GX7ĥ�X����4�C)��D3b������I\���@�[��+	M��A03��㼩�ݠM�g����ݲ6�j��jW)`�`�����'��8Is�^W�^nBc��0�x��/;�u��sea���kp�X��F�J�ՁGږ!{��<���T�<aե"��F:�H��ӑ�)���
�IJ�t=@%3��O�2���-�n�e
U��<j��<�Y)y���7�{!�:U�\�1�U��n�#gYE�\����� "��z9����Kg̯������ӱ��4������;d��Ke@Ȕ� �8��
�|s��u9�q$1}T�_T�uݯL���]����d�0C�~�m�}��:������RX���0D��^����r9�D�Y����E]Jd�B/�M�n�b䃛�jb~4�^:2H�*mn���@��x!،�>�8��K�S�C�S�Η���Kb�dͬ��Qɨ"��v�I�"\��_}�c���K�͝0���Ż�B���<r����X��l𷸸}&Kw6O�W%ʁ����ǥ6�]����0'ӟ�u��1�1�Z��-Z�H~�ݍrg��"T�:��a�u{�C�#�3�.��������0	��at6�\�r�eA��.�K�u%�0.<-��TF�����BS�H����.�d�K{{x�e{�綍TK9n�G�T1%�ȶ�.$5W��=�dt����tT?^O8��
�VO�,��rbJW�%�2�
� � tn`H^ $�.P��.ÌF�lH K�1:ӲX�jN�3W6[i8��pE�U��]�R���Wq�s���n&{�YH'f?��.�Y?>pQ �0vj���E1���WC�V�m�����s�8��=�p�`+mI]���G�R�����x��,�.5Chw�2`l)��S/g�v�S2��o�}(�˩pB��Y��t$|�{�6��/I�¸c����d�Ϸ=BjR��Ʈ�����q���&��1��Ɵ������]�c��~����K��G�d"��p�-�I�>닀R�e8~	d�-���g�B�<f~Ը��'mT���b��f`
�<����Jʝ*Šk��Խ���-nX�����9`�F}���.M�i��>:�<Z�(�Ӭ�J�7`<PI��lj[uE�.�W�'+`�Me,��â7,
��-m(��"���W0i$ڌ�p��mR�͌X�6���uvh�P,���&[{�b���8Y�`?p�#��P�T��gK2�Ϝ�E��j$ĵ���}L�K�ꍻz%�>���xqch�{\M����@?��b�K=��k�6�n&�Ig��
��T0��F�1-�XX�}��#��nFQL���@0��3u�'�ɩ^�Eڜg��j����R���iTج��y�:R=�t�?��GI�}�d����	�d�<����؛���E����')J-l�ȼC]P��&f��Cܙ�t«.���i��䈌��^�E��	[��9bMr�!��ף�����e��j�9���s(��W�	��0j�փ�1S�-�><kqn#�e�;œV��Uԓ����1�s��h"�ܡd�!��/2�
K�����8���i#������ v�~I�#��p�3��ak[�z` ��ML��qع��, jǑ'��]"lՁ��k
V�o� (�l����b�S�Z3���PQ���F�t5�㔋g2HE�?L9���~}`Ǭ1%�GuV�c�-/�-��\�w�29��$rzL��M��f�l��O1�jf�$���r;��1tK|	�ꏲ��RC��c�<�$�s!�f�!,�H�����m��:M�Ϛ���IpTn�����S��]�� мej1`�`tY�s��Wd���N'<7:U�Dne�ftec�(1�;nri#ܪp�Q����z���S慟�zP,�	x�O�_Cn}�is*kxx̗��~1�&��i/ĥ��Z��3�?�	wc��T��x"���V�Ƞ�c�m���C�U�Y��K��tw��=;�>�\����^
]6I��"^\���d�B8"�?�����y�8O!�8���%n�!��a�ފN��,���,��sCY#d\��A`��G+�x��.�	���hm���e���U8�kK��n�;�;���F�B�i	�b;C�y�6i7͋s߆=�)�� M�:���6���{�[��
h�I��@g<һEʢ�k��#Bͦ�x�@�C�,�`4�!��D]c�eV�/`zl�Jr`�2	81W��=ᜇa��	����xUY�ń{�x�x/�{F84צ�EH�x�OڳBd�A>s'e!XRpb��6<�
��W-�D[iS��l�t>�x=Mw��#;��ԝ5�����d:;Xې�H">eh�0)��r��0{��p�r�m�X�	��
�Z*�]6�ys�{�#G�pY<%�K��aC*�ߓ�L�n��ƵV��}.z�¯4��������o]Q�r�*'Ok�7|���/hI�-�Q�@,��G"�?�zR�����[��_��+U�ԟ'��B]�2��4���f��F7>�pC�6����b&�crCu���i�W�0ݛ����w����ϻ3"=Ņؔ �i� e�͒6�ZG�nC���\ݕt���I����F��X�4.���	k�O�"����� n*+1�d�S(6��>�2�؁�T��"�l;�a���g�0� �������{
���+ƶS*��޺���`G�4)e�G'ϛ��f��8G��g��12��Q.��f����mޒ��P�PYy�1\i�ວJ����{��Igk��y�s�����`���Nb��C%���&,ǙR*��q�A'��]T�,���m�s!����|��}��)��w�W�K�W�y���g����S����p4Pp!D�L�D@6�W:c74,�0���~R��Bૉ��04����hHk%�"9#�	��SI`+�r�=���J'����%#*[,<���i�VA���G��or=QU\UX|_LY�Ŧ�_��Q��Z���PΧ��g�+���#F?�H��a�W�x˚���W!�k��n��:o�l�'��YmSH��C�e�9���OJ���-P�x�sC�V�x��e:��ɓ��J̸S�#�5�Θ���f�����@�`��������G�%3&��%}ǀ)?�"�n�=ƹݘ�#1���o��Ɋ^qPY�^���D��%:0E|����+�a��J������Օ�^��W�E�M歞��r�U/�� +������8����4Js
��x�yu���d�B`ax<�]ϖ�e��ƒ�)e���oc+�$2��-f�`E��[E�.r1n4ͪm)�ł��0�&��� I�؁(�X��`�ze[��ɟd{ rkNJ�E(�a�h� z�Ivp~�S����QJ��w��&M�k���Ő`Hz�;x��cYS�� �ؿ
F��u����>F^�c����}���nQ��c�(r���HV���6��w�|�4`����.H�aԭ �W�ͥt��ƿ��p��V?)��e�����3�ьIS�f
G���o����t:5�&�Z:�g�wܬ��C�ҙ��.�/�cX�(�})6�1��B{{���Hw��7�~�u�a�j'��TF��xb���?T:��S������hRxG۩�[��A*)�[��_P��U\�������>��H:��(��}T�zs�2�5+Y����t(������
���p|D��y�t�D�O��+�����h�
��j�i�f��8Mi��^nT������2�x��D�B粶(d`el�SV�����8����`��;@\:IO�lO�6��*uM�i�Y�شHdu���-W��ܕ����^��f`�+����`�z-�_?��ͺ�Q���P~�HW5�Yx�� ~����ʓ�C�L�C��Ǒ�h�s�UE�Q7
�f�HY�u�9<Ω%%x�e�Յ7)I�Ĕ��]���g�����1��,�*ʛ�>��l-;R�$S���K���:%3�ފ鄃`a�C�"\�n;�-<G�Y�XT܇)�a��?��V� ���#Fqu�d��ǋǛ.���Lf�rq���ޏ�!UZ�~��'�&���P^�����E�vJ��T`��*Ɲ���V�=cQx�GQ�R1W+��Vڞ�[������a����`����a3��ׄ��C$������ �|��Yf�I�g%/,����z�F9'�Kz�RSW�����N%�����`�M<ᬜ4�H\-��h^z.�^;׵�u0��٥�[a�Ǝ�ts�R�X"]���䍞���	]�Z�K��
�E��ڤ?/�u����!�:
�g�������3qnX)�/'#.�)�O���L��T�xB��fS�?>"d0IV�i����u%kB%���ė��:΋dl��l��z^0䅶H/J��.��o>I_�Pi@��Jv1`�.#�M��n�?��ih�5�iD���>O�[>����$��6.	�*��!b�KJ��E!g���U��3u�7�3t�T�瘠Q�M}��n<��cXΚ�n��/	J�ۛ��h�����4����_�Zc�>��V���G�*&A�^
�����2��)�Zj���\NA�GJ2ߴm0(����
�v��D{�ʢdy�C�@��N�����\mNq�8i�iP��Z#>��j���?�w��[eU{:�{b3W��`Uu��ދ��@�>?/u���;z1%��`��uF���X��^czOi�#o�"�W�*Ղ�3��p���'r����8�Gr�#�39����	d�k��1mVdT#��g�cH� ���� ��(H~Ѱ$O�{��t�y�+����� 6��wL7�uZ��Oȑ^>+�����L:+�����-������;K��_;���텆`�?{��%��-��SS�r�����b5$�!� ƺ��5���e0%�P	��,j7 zl�0@%=��8k،|칵���;�y�^����sGoۗN��M�"�٫�􏞍���z�6���jҠ���j���X�#'zt��N�]��Fm�'���U�|��`�K�����q��*,R�
��OI{�����
�N>B�����ZY�"kB�/w��՜��i"U�[#���]h>�QѸqYr�&綷��Mu�o�c�7���N#A�{𞐙��`6RGEa=&� ��H��SO�}Ƚ���i}u��9¿���D���	)�NJ{;�܀+�NF�9��W��q�ߙ���M%���]�]C�\+ޗ��K�?^��cb���7w�^:��+D�rHj;�!Q*�b ���,ʳ1B��YO1�8X��?ݬ�>�
��P���F���w��sʴ�Sd���$0��d��:'�:Tnf{;�u���S��j%[j<��"j�ʠU�vKR@Y�R��\�>�i�D�wR���h�3��jpn�?/�
��M�wǥ!Q�H`��^�~+j]R��ɌH���X�eY9�:��-�H��/>d�Qh�J"m.[���"-����1R��	�����x�K�\�z���o�[�3�Nyۄ�cg�A\�,���:z�Qw:���;��%kc��w�0�Z�.���y�qYm�t�1) �-�1 �lk���i
������X�������U����`�9l,�;+	�wg����=_�k�ݛ��f��1�M��h�N}��=�g���\�Qx��fLe�29ui�����颠��YFy���CeV���'`9 {�n�W����	ʭ���~�����t�?>|&0o�E���Qn
�-��(S� ��h����W�t�5�(;��Y�F�z
�*(�	�X_��7ZCx���5Ś�@%�&f$+f����}Lκ��b�9,{ئ��]����oG��,R}���%�(�@���,�l"mc��bN��`��+�Bҭ;���e?*������ �FT1 ��4�j�TR+���ye�[^YFCA��dj0CfF�q��Z#�V����t�\��$���>e���-7��rXj�wu�J�)Q��:<C��j�{��rI��2pGX]�(W-�$V�AT�K���n
@�A���m9��X��^[/���s�툎c1�e��$c<�B/ѣ��&�TI;B��LbҺ����B��)��˿���,�5�����vI������p����a�@Q�w]�,�?�k�g7��)�B*v���?e��lO���SY���+G�03��(x�s��z���cGYGE����RJ�2�iqQ�½?sM�r�_���Şz�d :˵�Yh̴u��;[A<>û�ϫ�Ek*���sŽ�J�&Q��5ȧ��B)�~�o4���S�]�Q���Uo-�g��[�F�M���l���D�X�� ���5��]b�uF������P�|�Ql:�m1�Bp+�Wҝ%�s���6�_�X��7�n���������*50��X�>o{�T��뭆���'�)�Y����w�I䴰�
0�"�`�j~�|�a$�16Z�N.MF�}M.E��+�[#c =�{��Ͼ�t��G�ѫ���m���O�?aK��In� �$��>y��=�	���F��Җ��U����!��3^E�,���uh\����_�k�� ��i�  �;�����q��#S��+SS�"U��@G=����%@v��j�Ki�uT%.s�G�H�@��s�?��n�^�'�p͎T='K�5�W��`_c�<!��
�m=�}��U�bu'�"�h����R�!�a�Ԋ=�3�`Ly�iF3���W�xֺL�+��ڑd�dNǶAXGn�Y������i=烝8��q}��rj�'~��#�K5t�gu;T�8��֑�%C��_)�Q�����Ux�cl�lV��?"�~���̜�E�uK����X���nE8^���TP�ᬗa��N0�����8�UA��H%}��0�7b���ہtOa�}�o����c��i��c�|��4Λ��t��)6��%e�l�}߉�FB��P/����y��FwLX��Z���
�����W��&l�pK����v|͜HƄs�l��fԖ%�б�;:f�ָ�޴���b�55�	tv�Y�Q�#%��T*L�P��]�w�yhG�;�X���	�0�����IaD^@�V��sڢ#���G�D�.![iQ�ك��c���=c����w�L7n?�k�5��lI-S�����@��wѲ��{wfI�ov�W����6J�I�A�*=l��KūK���Su(q�{�<v�U��9��(��'��q�f�V��E�u�2�ޭ����A|y������[l�R��p��z�|�Y���q�����:��?z��<�������ȕxbf�[n�8�8EJl�˨\�	�5#�}q�BW���2���g�a�|��&��O���V��#��. (>�ld�.-e��������7d�PC	��"͔*�^1����t�{P[�����HѫN�*�sq���H�
���m4���$#�[.�A]�:��l�Ky{g�8�V��j��I�u����y��tշ��1���~F>?M�oJFy+��w��t8$b�{U砄��ͣ���h�c�Ux`�P�Ǣ8�O�����i��r0�P0O�ڙ;�&�"Q1�
w�����t��Mk�Cb/
X��~z�Q'=��Y�ᔭq�6��*�~��@�Uw- ��M�h�^mܵ�}bh9���1��	�2œ��\!�����:�i��0����x�� �2ԖW��[�cXv�.,��f{.Q�����6D��|����d_�D#�$1�0/�شk�!3��q�R�������<h��,�T�F*�V�S��*x:?�F}�}�K�#��܏f��!1?!̛��R��ڦ�����v���K�ɦT3VېKm���!jݣ[��
lӏ%���t>N��+в�K�d�`\O]e\剠u�(P=��%f۽������^�R������mG���@��.>����L0��ý���$�:��]?�������a���dc?~�%���rd��y��V�W���v�=���D4�`W�]�M�41:��k&���.$g5\���_&����B��T�c�#�:�m�Uq�;�4���<SR�G'e��*��hp̅z������� 6*�6(��GF��C5Q0�8A�ǦaT{���݂O���7q�/.��������%f��v4�A�K�F�J?J Ypags5����`�g�)�3����8Li
��amilW]Q���E�0̿�=,O��&Vt=��gx�@*���v�\m6�.`���� :��b�S�E$�R���˚RI~A?�b΄��	�;�������A�����*_�4n����J�N��@c���!�Q\d��3fG̤�y�ݵ���u
�X���g5#T���"� ?weB�G:�z��J�m7f_S�.{����ʎ=3Sډ#���,(i1�a�;�hj��E���� *^�ٳ�5ڪ+�Á��)�����	�|��6�Q�$,p�-�C�����#�"&r�~%�}Fm�a�������ܻ����r�M��!�|�ʯ���r���d3��}���B���
<���P+�_�Q���s`1��)�<G$l^G$�����w�M���j���]�m��O���SlR�b��� �f(����
��C�I
�J���Ձt	�U���[IfY��S�l&4����~OZ%��2��l�`�i�*������ԋϠ¬�hC,>	)�J�F�����'ږ�G��"�߃��6�WA�f�Ǆ�j�P���E1�����J'qS�ק�+Y�����k����}��_�R�W�1hwW;_��!:ZK���8*�?�z�C����eR�[ɚ���05�R���%��}�[X@��ċr��Ҋ/����B%Հ�ܗ�|���(���u�ؓ��0����*�Ө�,���^� 9�����g�L:�0,V�ؠ�2mS�-����R�q�_L������[�&���2���8�q�mGo�zRytgb�����@Q�9��j��'_H�tW��	i����O���̹�ۀG~HJ8P�_o�9����g�OX���yϗ�JJ��zO�}" ��}��jK��:Pa�)�^�Q��9��%�ΆBTzO ��,Qf��ec
/���`�{~gyi6�]��1���I�����c^/&�,���
X2�
ٯ�V���i����;'�cʪSN�ܘ�e����0�L`d�D������>i���(��W0�t*r��>�ծ�_��m���m���;��9U��d��T:R��oOZ��Y����t�뇉����tI����7�	�l/<шL�ʔ�K�BT�ag$JL��Nya��x���Հ綆:Ĕ4�݄q�!��8'z�����h��Bg	n�R�Y�E
~|I����b�!��=�3f���[�<b�V�欞Q#���BH��ҋS����,��A1a x,�^a;�W�ǵk����L���MWj�|<�ky8����#r�x���I��%�hj����d�>�J v|���ML�^��2x���Z�~���o,�ʤ��9�	Pa�j�	q*�ډ=@�T5DSX��7i�sxZ��\�G��!jӍ��
u�
�l�R�ѱ�P�Wʈ��=�yQUy�޽^��.!"�J03~�S���'���TS�$�^�@�(�h@�m=ltˁ^p�s������ۛ�QP���� .��.�x3��ىn�d��Y�]z��|��m=��vJ�Us@�o�EL�%���DՓ$���E��I{�U�2�ߤcE��
r$��D�2ٟ��n;.Tg�"��^?r�rt��L7��4J�b ι3ٓ6�e#��-0��p)q�K��U[��b����?��Mix��t	�l�\�B���G���L�%��p#�>�S�%D�o��n��	I����bmYA7�7��hʭ�1܇����{�콴�m\����a�Kذi�ć|
�@u��������t�4�S����*V�<��o��|�yS���є%�kX�8Oպ}@�v�>�Dq�I��@�#��˰�8.�L�͛">�|x���hh����+ŋ�ub�����5���N{d���0j	��+nM���V�siVY�YLm~������,�5H���cwn9S���l�~����	�>u���!��#��߲/�X�r�I��{)��0���p�f��I��	��\j�0�x����p6�ǐEa��n���F_XZ�� 'JzN��g��{����j��E
1��c#�҄/�\� Ҷ^ЇE���C���=�gN6����^���GA���O���"哉�r=������/].p���ϟń@�vկ�,x��A�_ܦ�|�=�u����
I���^�w}[,� {m�8c>����#��oV(s^�A��fO,g�iG6?�����MYS�Kqy�L_���Bǲ�E974������Z8:W�˥�<��>���JQ�ro���J�˙��^�1:|eW�#�33�u�(�TG7{�j�cwm6����W>;V�F-zds��B���c�jf���D)tg!�|�I*<��S�-@:�2J��Ъ�uQI�������5����<�(����D�L,{��B��1.Kᛴ;��ox|�[��#
CA-2s�,:���� â@Q+h�ox���=��%㐶H��m��Kz���yp�O��~㢉p�����K��Z��ʃ�yƦw�wd�*�!G��A�M4� �y�=d:�xF���٩�~L���_��U�忞N���?�g��
{�$��������r����K�QC=�ʂu��^�_�r��ک]Ťste�Q��7GL�����������f�26���%1<�P)���U�%��C���s)oT�����9�ij��~b�_�UsS����<-o8P�#CO`�����@�aiB9�	�<D�Q ���Пl�C��e(�ۃ���3-]A��Jh�^B�?��'E�
�-�vXE�0�3\ߎ����}|*�7B�>	����,�;�~�w�+θΏ�͒�2�J���˃l
��9��L~��@P6W׽��b۫`�kO��W��B�|+�]	-魔>5�l����zۉP���Ը����Z�53{2��Kã�k��M�0{�h{���%SkA�E�(�\<�cz}��1lߝ��SuT��$񚫒Z�N��g57"lNu���y�<_\չ�Հ��4����qY�d�{���	`���<�i�&r��x�����O������e֐^ �8bةW���v|>��/�H��8�l�y	N��p����xu�N���aE�Za�_<��k'��lM
�d;*⒨^d!Xw��m���c�;�������7�u�l�~�`��b�T���h�ӟ�foQ��$Pt4{2��̉�<Y(�L-�YR�ώ�M��q�FwH��CG��A'K���7g�dof�q�g�\N������r�V[vxa-}�R����n���������-n`�oj:8����KͰ�2�avYB�](4�㲖�]R�M��3�:�t
��	��
�����G�4ܰ��¢1_�x��EGDk>��p�",n�m�?`�E��ͧ.���<�_��7n����؟�`�K<��m.Я>��F^Sok�3��iՐMF�.y�����Q:�S��/?42V
�|D���`�vv+{��M��{��@��F���W�RN1�W0'�
\�����8F�m�$��u��nmj	6�Sd��Z��qe�Qnb{vn�������hPJ�s�e���1i'�@�N�D��ԏ
��V8U��8�čI���DI㌖f�2Wgb�*W��J�!{��肤��3�5�:���f�מ�5d|8���TX�����R�I���T���>7�>!#pb0���EdE�M��#u�>��& �=����֐���$�j��[�6܈�Y�	g[dZ"YsP,��	����gP��yK�����mϒJ�9��H�9��;B.cA�!�����3\m��Oz���Z\ r��?
KحC8"��>Җk�@�26=��_0���(L��o����I9{���٘ܫnDY�|@��8jTF�����6*�~J`]������	�A�u�~ؼ�4����/-��������Yͽ����ٔJ6��k�pc�R��Z�w8u����ѸyM�s�@�Q#�k��5%�E��X��Oϻ��A������?@��}W��:�uÖ�KG�
\.�^�3�Дg�p[��d�8V:g�Hp�My�%��#���A۳����G|��`Y"�2�C�f;V�kH��|�k1�Ր�����K�( ���bn�����>�o����a6y�}���I~�q�1�� -�M�H�n#x����nOI�xN<���^;�jȨ�9�Q�׃\��[�|Nm��0vA�?����y��y5�h�P�l��7�+!��2>@Φ[T�O�D|N5��[n��w<\��b0��0O͉V�LPӂJ�q�B��5�F�������O<��C#��N�@�]�

��G��Q��Ӏ�3��fY/p����ⶔoد�~�-� �A�������#i�I��Fzt˭�[��;��\g���C����]~����.g��H6�r�s!�b5��wp���}�N:T�zߓ��|��%,�^���$%Xenm�#�3r�b�M�Mk�E8�r&�,)qr[�T�	���#Q+@��0N�\�);��oj�)38A���<�/���o�����ӏO�KT�Cy�O�>�mP Qu	�l�Y��#K4�Bޮ�ڭ�fAM���3Lg���������O�p[$��mi�
��2�u�MH ���>�Sп:SI-�ؘ�fta�tz&L4k9����3�p>���������J�f���B�RX�˼	�6f��ĎajDn`,��h�'̺��lh�[3��}�ef������	Vj4�"�E����=��eb���\�nZC���B�*���@�w>� ��z�Ӵ`��&s��ͯL-������RA���A�&ь���U�e9�'�x�o�ν	UPD��'(���,�E���s��[�h#�v�j���Ea��.��W~�~�I�1�U�����g� ඥ���[�O���ai�L'>0�d���0pH2�{0)ǯ*2�]���<17��맦:26�����L��s�q��7��=P�{G�/x�J��{���)n ���K&��4m)e�o�ݧ�����m����M����2��{S:}����@�..CWX���gwߟĖ3�tD��~����e�֐:&f���G�38���$a�D��籩�QĽ3S�\�r�V�Q-(�J������p�.��E��(�Z����4鋦V��i~/�X!�7�$c��+�:�kz_u���3\��gJB�x��6V���R��p��G���e).&�_]�������Z���ԗ94�1�X����4��B�F:����#?#Z�RN���<�V�%%�����SH��z�I�qRU�u�d�'+���O-�H�X��%���8rcS�e�q�(d��;D����`�)��n�Yd�K�7�=�I��2{0A���Y�o	�Q��������5��E�	����������4n<M�;h��#T� ���$&������tm@��f��K��0���Cc�MH�!0�����w�x�� ��g[#'{3�J����s������]�e��������3�E�bN����N�_~M�`T���L1>�v�Ȼ�d���"�l�9/5 �藬Wka���*#���M~����p/�7ֻ0���u�@�q�n��n�4[��2&��e�4TC�����^�γ�6w���������� m0uID�=Y��M�>(@�:�^��E���JhP4��g7�(�7��h��o��r�P��d�*%&��.=�Z��T��Ad`�	J�����C�ڭ����T�S#�D��$���8���	���N�I�+Χg#gƴ��D�T�e��Njq>v��0z+�(<�C�����,�^�1Y�%Yl�8�X{�i�4���;Z2 �����Ǧ�~��J��K�Q�.���iJk�3Mī�jf��U}S�8��>��1xz��lSܬ�4�D��[E���<b�����5Л�.��'k�r�2Q�I�Šߋ�o��]g%~�a�b#)�~��:��."ނ����8�G�[���	�sw��]�y����ڐ
���u�X�սL3���o}K
�H9��?�g8T�h:@�xbQ�������v��C]p��� ��#�r��_?�t'�ûn59�R��E� �����7DJ��Z����G�s�U�v�Uݧ�Ҩ�_��01�5	kv���n�@k�5�$�\�_6��5ⴇ�a�\f�d��ҋ�PJ �؋��G��uN����02�)�kõ��%�K�J��Z�\�]�j�l"H�f&��>.�
�"I��[�y�%F�q��S��,�P�eK�;��\�*�jD��}Z�Z��C)��5Š�f�`���P'���y�P�h�<�='T��B�GiGp,���51��AJ�z��L�d�%���������HFh��˻�o�9�d���J����K��h�����o��^/�O���a�GțG��^�"ɫH��?�f��rh5�@\�\i��S��w6�B(�X63vv��#M��c��6Q��eFn�ܨ�+��l�����������'	�J~�QEY5G�C��'Q����r�!Oͦ���T�HM9̾�QI�5��+���c!#@�h;H_^��iV�Lݢ���2)� �6F	h��d
�O�4(;�<ON�ۓZ�4��y��S8�Ui��s'g���fDt?dA�C�9[U�#o��dKq�W��"��븪���\�#��)�OdC=�0 j@8!��$�U	���#�F�3 �1�l<}�"��>�O���e�!y@�ن+s���X�p)��A�ń+1���H�ow��������m����k]ܸ��O�TY.Dz*��01?��|2��Q7\G�M��L����ʸ� =�d�1�PFQL���.��qr6-;�[����Ed�Ȓ�%0�f��L�����D���ڽ��X(�4a0t��w���A~^S)��8�%l]z�v���'C�������-�{M�U%fZB�,3\[emX�m��R�e_!8�݂� խ6�qu��-]�!���`�1d/I4dV(��,�2yC����޿] �#�1,im�$ل���G�*oI�ZHe����*�܎��FAC�EL�)���!�	�h���2���U(M���;>1����z�O�V�4��U�c8�} ^ʅ� �^����h�ˇHO�����#�5� ���_/B׵:�p�f�"]ޮ0^%IB[4�zft�he��Ӵ��D���>Ռ�]9c={݊�#H��L�_c�tO�ӧϗ߿ڥ��m[`��93�E�`U���,�ePR#Ad�u@���n�Օ�(�Frw��̓���ha]���~g�/]�)ɑ-8C�Z)�G�&'<`x:�!d���96y�8Q(\�ʌ���2�]�ZVj��ʊp&��]�ZGG�?�@��?� r�m#Q�`�:��_��l7���;`��CA�k�P�#g��AU��z8�Nk~�� Ю������D���W~2��t��L��Of��?>�2n��$�-���V�����4&ÿ��nxx8Ø8�V�z������t��Q��Vd���i/�g��YF� )����- ;L��9O�+�@��B��0Yȥ�t�-F�\�ڷ[�#lVZ���aĖG�fL�z��ֹ.
��ǅ�s�Cu��,��h�Lr���e��Dnco#���R�33������4\s�,�Q�ʗ����w��v�uRǋE��Z�OE_{�Ȓ=w$�c?���	j��T��g!GI����e�:�hL��
r.u��_<���5R�d"OK��|oOe�QC�sͩ�3�h�}��{��拜80��*��G�V�E�_�Y�9�!���+�W�x��K�!�]��N��w�Blٓӕ���ϩ����;7�>�4� �It��Fz���{�~B'���I�-���H� �`2�b�nAԭxw6�3DS�Y�i<�)r���}�7m�m]�C��O�0��5�a��v���%�ĵV� .E�K� �we����f�S0`�'�o��tD���n廄�;��E1j� c�u�r�&9���c��J��h]r^�Ttε��G�����m��l?o� B���AR�a�@��G"@+�6�4%��!K��˼�y,�(3��uZ��
%�����vf�����&2ա@]��ޒ8�XC����w�Q�X˦��ct|��;E�K��aĳ�Sӆp�^���c@�����U>!�כ��v����l�W9uz�$7a[4��3�Gܖ���o �B�� �fq��s��3�6�k 6��]�����t�V�Ӳ	�����.IѢ�Pzǹ�t�h�{q��wj�7��X�������W�ȁ6~���χ���q3.Z8�y�B�9�H��B%e�V�~�^�}%ǃ��N��w�2��a��W�c���'��9�����#�\�1�Վ�k�5��_9��y5A��¶S:�$	��-�$�~נ3c���Җ!�k���@T	��OJT���L��F#'��4H��k�g�y0�H���.qH܍���e|yL6�lcb�6���D�qB��푭���OY�*��;��@�۠m��M����ߣ>�7o�y����ߡ�7(�̻\����[��&�td��k����F��-��j��ln�����'�cm�'�+����|���e�o���	^�����m��,7�{�e�X7�iDI�1��dB`0�ўq�c������Ul�Zb��m��R���y۶ϽI���QӑChJ�q
dC`�{�9Eg�SI㉑u0V�����:�
\�/�>���EHEa��߇��K����q�Jv����E��0/���N����g�
�S�*�BI�Vi��x�Ɓ�k�6��f
�n�L�U��O����{�ZO�0|�|�I��+��uT���F�gr60eY^��v�����7��Q��|Y��&�����������p߷dA�i�j}�9))����=�U0w�lY������C�٦�?N(�LP�5U���w�NE��"q����3M���"�gCR�(��D��w'�T��w���j'vS�4BW�e �U[�/c�p�D����oa2����6�����ѕ��dq�����]�(풤:��+ey�L�^�v���2�r/��
�(�	)	�V��;���6�;��F9��
R{JL���`4���*6Z�C:\�8�	D�	�)������o�	��7�ן����[f-|d1:N&�&&�z�����b����F	�:2N��(�*�m�����Ȩe�~�H:�0��)�t��b�0�p�z��^f��@��?ʹL�;�j�O�*�K^B��e��G�W���ߔ�Ѷ��C����{�
z1D�Ǝ�̳A����2đF����M>�=��h.K��m]EZ�ߑ�jji���s?RK=D/۞���D�B �����F�7K��j鮐��g�	=�:�A#qٍ��S��KkT��87�{{�w2��,#V#V9�a� ���z͐?���4��?v��-z"��Ψ�x�1u���$م<��x�S3W��slAmO�v;u�"��iB3}�ZaؐU��a��=œ�䃦i�]kt������b���-R9�8���t7����'�	������761q9Y\�X[Ā�6�L�e���}#SF�G��E�)�w�W?Tݍ�\�bf굍�e?��+�Q��b��Fm_J'Bs 5���g!�N
�~��.0ПaPڱ������q�Cڧ��G3
Z����J��Z�~�(�.����ă_�`�����6��5n���U�p3�Ҩ���)]��F�{����Ij�־��~9%R��z26��A�N'�W��&����=��[�/ b�uɿ����Ԛ��d�@����� ơE�	��^`nj1���טgyPHD%�D��V�T�'� ��(�>��9��x'k����Q8y^�*n���O]9��2��;-�:~��3д�>8�I��'c�� �PƦeiޓ����c�w0q���k����§(_�9�ܸ���޳� $�g�P ��U<�#1|Xٓ�]��@���mN3AL9d\�p�@G�b�����A�x%G�W�6��s�ZjI�E�muP��ю_�=��:&����3��ʾ�%��/�:��U�����~�$V�f��� ��(��3�y$>O��t��fi���GF�	�G��N���-s���'�W� *�2��� ��O�8�W���=����w~����|���p�Ǹb���s;��Bx��kWׂ�#s�t���Y��`��?�(ő<��2),_�\�DB�@b����4���<cH1��3��~p1j|뿖;�mQ��鐢��~qҺ2��s�W�s�ɸ�Ek�1�S�J_�'!&��'	��i
u��"O�S>5��X�$m���Ä�gⱤlHv���.�,�5B��L`�|\�oܖ��8��X�QB��ȠKKD	C��j�%$���,�S���Ø�}�hB�Kނ$O��L�M��g{n�y��3���yn��Ş蛽���"g_ ª����g�ʿ�{�*c}8��O����hJ[[u�һ?q��/�N���["�yX�o#��8�Up�'Y��[@J�U�:�Vw[����BOn�w�:�:}�)��F5��تy��2|hs\��"&���*#w�Z��CL+P��e�O�}�_��?��G�I��/LiCQ��FF�����E�����b��<ߙ�ʗ0�ŬŬ�LM�cm�儼,-q*���3��t
��b������*�:������<�z:X0�m�������me��_��!�u�pDV�IZ&6�B�%K����Z	 �t�A�?��m�O��r��9&o�+] �<J�^���Oݪ�G��v�Q�{Gr'#}!�<,j-��j�ކuԉL���R���я���_�(G��g�-��I;�7�1#����b%�KX��9��E3���!ҁ>\��XS�1��A�cꇉ*��7���������O�d������1ϯeuE��2�J�����0 ̢�P��:�f<|L�E�PX�g6�5|�F�fI��s��<�+���F��p�j@��pzF��~ʩ6'm���`�x����_�"�~4�4{ <ٯ���Qx [&)G`��M����˘N��X�@�<��t<��=Cy��]�����u�������
I\�<�F\|�w�;*��<�p�Bh�/+!)Ğ�MDo��kɋ�},x��"�Ig�YR����g�ic�����a�;V���o�6#C���(�\�s��3p�Emr�`e��;���ʃv!G�I�W�n�$+U�� �����D��h������QݴA��M����i3>1�U��L$��/P��0ӭ��>�ҝ��m㋙l�ɋ��UR����<]>+���\�j<�k��	jab�P�[m�
y�aiML=�^��6�=���%=��
GG���Q������0�xr	��~(�#����sF��^���fU�8:�bv~�d�U6ϥ�f����QL�|Z�$V�6��
����*6s�eO�%gd�����0�G�d�f@V؝Vn9q��G�Ru�}�3���AK!q�
�)-P��V� Kf�w�le�+�{�0(���,�i����?�B*b��jp�;�*�k���ta��*��ӕ,۠��Y
[\p�<�-r��'Bh�a���ԏ{ʼ4/��p�}9��^7�<��uͮ���[T*
C����}��Ș�1�}u�0�O۾Ny�H�K7�=P�Ntd2�g�ӕ|�;�4�,��%F;���8Sh��"���`:|�q���6�� F˻�C�F�2�������8m�B���g�8���?7�*�S&��-W��B��tJ^�W��m�?\�+�>���cو�#�V�B������/6ӷY`|�x#�3<<(���(�Mu'>k�J\%.i�g�DmQ&ɦR�R]6U��ѱo�ܷRf�RaÀ�?���]Hz�޸�̴��}�vp� t�l�(���<<]P5��8'���
F�����6���\rN2���)�<,�<����仮�~@��TF5�������؞�3P�Ǹ��w��ǅm��.xp�n\�ڵx=.������ �F����l|�w&)r�ćE6Ǣ�Sbp�|{��n�,
C��$g��D�+Iv�3��!�������de��m�޹]������*�V����p�^`ox��:��US�\�z�ʛ|}�)��/�v J9��3�G����k�l�j��$�g=ܡp"�l�yS���L�q�n�a"?����M	��;㕺����P��`�PW�c�-��5�
I����*'C����Fz�� MS�i"C�Y$a��k�f�g��~t$������c�}^�N��u��_r0x�5���Z.��+�BQ@LU�E���v��F�>nj�_S�LvX�g( ! �ֵj�0#p�$�pg�'Bl~�uh�l[���$ �v���>BH��!��_Y�'ðϠ)nx
��(Մ�/��;�˴�xU�ɐDJ���VRB���$�hvH��.�����B�B� �e�r2�+�@��o��mH��rk9����T�V>����D�bzk~Q�H�Wݙ�Ps�ñ|�o����eØ��������U�Gd<�gtVO��nt!|�B�o~)������+`��"�qI0��lt���=�<W
dvzzp���h��M�������a%�a�k",!����V#��N'��s8//G�:�3̦��KD6��tD�����r���G;���7����SH��s �'�q� �w�xcVkD�Sp��c���ߑ�Ѩ�տ�
��Aj����pW6@K�@2NB�E��6b�;֗�8\�6babYX$˒B��Ʀ��+�#k{����R�;�w� �r��q�(�5U����~72�72�U�c�@sNW���00"(h3����*��Q�5��(XjG�<
T,Kg�9Ԣ����R7&z��=� NjO]��$�ԅp�>6ӔEb�����;Ӷ�:�V̘�*�3Q�a`#×�te���*'�]���	o*��b�e�-���ysy�z�y��s�G��*=�u�x�gw�Os*��[��6��Kڒ�5�R�m��?A��Fz.[q�=r�u��s��%�:Ɣкkթ=Y.^���F��y�#�8L{"�>����e�C���Y�M{�/'x�KF�О$xMuR�.���ϣ^"�HL'���4t�6���l�[�VN�i��KA<���o�Ҿ�;yvr4f�+>
8�P��ÿ$
z���|#��^��gL�T�T�	�^!�K�fTO�ݬ���ol7�,C�{:�mb�V���a��hK(� N�T�q�L��נ~%J�r��cC�p��<�Gs�[(*3j��B�q�^~,g�(.��ؚV���{��q-�u���L�i��?L)h6��]Ç���Ԧ���%�nm"G���n���o����?��W�KQ��ĭy��D�R�m�6Y�fvGG���0ZƵ���0��!��WC&jj�츰�%�#&i�:�7&��=5�]����Z ��� B���Z�5`�w����2Rȿrމ�q4�Pe���ʾ}��%�6o�N��.b��0uȏ� �=e�X]D�-1<f�����ܠ��5����(�#v2b+Fˮ_@�C�àGRM��� ��$`?b��kA,��c,�A�\��A�#�H+��?�@a�b�io�FPG.z�٧���浦�0C7�hؼP����c��W�y��M�Y��:R�j��cLAD
���꟦Hk°����?�a\��++[2�������\�l�X�X�rf��q)k�3-����� &��nb�y�2GR?I�g���R��kv���,�lb�ؖD��\Wl��,�F��R��Z]m6Ӂ�JNp<g�In9�ޕb ���.�E����Y&E�\�_Z���u�����<�}D��BI�oMx�p ��/�l�(���"�Efu��7�\�0]L�'�m$7��}�ۭ7)	�\[!\�����#����2���Q�oxTb�4�mU��)��h>=9k� $u[�F�^���8>L$nn6��I`���z	ײᕿ�(��۷FG��6�����ǽ�gv�v l���F=^�0�w!Y��H�#X�a��z��,�|7�f�L�I���<s5RI�+^����ڇO"�>ڲt;<�s)d���8O+��'���"5�뇂/�ř$-���[v�����������x�;��%bs�Y���.�w.E�M���v���|芖jS��Q�(
��Kc�s�7��&��Փ��߃ի�V8RP/��_�ܡ^>��O	����(Z�� �Du�.�a �Z�*�0��|��
�2�X�%��E3�l�R$y���������[�꼃K⏒	����bͶ��CZp�fB�T��/ T2x�/wu�BW�=�J�,�Pn��<xI���u|�|M�j��\����{���+�����#�$�'���&w����-�!=��y���
	��8���_�O�κ.��$Ι��{��"{Zfn����Q[M�D�4�8�)z�v\�KBVlA���%���P��P�`rL��9�u���V���L���Uv{l�Ͷc9���,&���(łY�u�a���ғj�Meb�{�D�i�&����ke��N�L��ؖ�s�G
:�<}��6�)��jOǔK��i�<��Q�C���⋀��oo�Uk/W_u�L���Xwa�'F@�l7�I��.װ��C�-�q"4"L/�-���H�����ƈ9"	�x��UL���s�����Lf(��DΎ��Qշ,,��4𠺭a����b�Zqm����S�c ³"J:���h����4�ؗ����;�K��oh�VO�DT��/Y��.I��}�u�����U�@|�,��|e��7�^��O��QFCLc%�u��!M���[�{!1�_8�1�C�a�r+�1��C�2-Is$�رF�U7����B�X�@9�l�0�'Z#��E#��P��4V���e6v���~��zym��AXs�D-�(؎�v��V���v���t0 ��BqD]Igg��<A�P���<�y>V;��U��`F ��Z,�H��ve��(1H@P�������O:�����+�G&�o'�X7�|D4ے�]�ID��g�gx|Mw��xt '/=�@�J�����0�������N����&��5��l��;�^�{S)`�v��a�6��W6�dS�^S� �����٨<=D�s� ���Yl����ֱņv],��<:2���MJ~����87UF^/������P�7<ӄ�=�>���@`�v�G�ě٭�֭��=f��ӗ�r�~3̢b!��⥰J��
�:^0Q%�d����o��C�����,t~��V��SbT]��v�^m�wEa���m��F,q���v��u6�fA/�G�6D���M+�D��@ގ\�p�t0*�z�M��UK���>m��zU|�~�܋5�䐵�v)�&~�_�2�~M�0��iB�M�<�������zKIɘ�'��Η�h�+��o;�lv�sn`�s��`���i��j�%ϫ�rD3�pG��l��9�'��7f-�&S�._��L�^.CB��p�I�R��Þ�x�&�tրR��=��0���%�����+.�N1�q-/L��yN�L�\�+��ttVK�H��Н[�* 6�wiY����?3�Y�H������Q��nJ���!8�I�����zQt�E�
!~���'�sHP;�]p[�e;�2�\�dW;f�9��8�{�+�0�ˬMl@��>ОQ�J`wb�2?���I�]xA��zϾ-�R�"Z`ţ�tp���Q������˨�h������
� N������Q�h����G=�⥡��{�9�\(l�����v0�v���x53H��m�'w2"I)6|vҤw�L�n�6X>|T~_=�k��.#:(}˓!~;�����>	Q(�>KTU�����#,�l#G�c�u�8k�W5��S�0	0�S��u��'B��B�gru��
=��N��P�FCB,�愌�o8�����L�#��<	;�e��<Q;+s��AE\��+��<`Vm#O_��&w�V�7FqY�q�ᚆ���#n�<VS�71t�"�1'�ʊI�� j�ɣ��t�xۄ�,�� {��ES/׀[�h����PH���Bu�O�cRHM���Ě�X/T��@af�@���Y�i����x����5,��>+D3�>�՛3�b���^yï�I��#���Cy`�b�eO�|"ր�A.+AOF�RB��C����5��^�o%=?ҽG/k�2Sc"�>'��&��9!�v���?��i2�f~ʄ�4����2	6d�It�U}P��x4��Ї�+�'"�������%2f`"�d[�AAW��7��x�#�|]�ͭa��pmz��A�#�������rҍ��{�!��v+���#>��v��L�~�]k������Ϭ�j�$¾�7�8k�!��;�z�(w��n�CS8FZT��q�f٠��8�L6�b2��J��uV�Hג�w_����Rt$T4*���A�����;���$�H���o=�6�+�Y큉����K�b!< )T~���v>�S���V���$�
H�.ѫ�[x����	Z)�Nm?�
]) 2��e�����1�s��d<8�t��l���9��g�r ���p ����&���[gGٖN����%�[����r� �t���'�v<$�j�PF�^"��g���U� ����ϭ��䯅�(A��W�&^%���80"PP�����y�m�N�=ɌR��-a�!�y�o[�����Rۊ9�sS�r�iʨ�pk���Ł�T.N��-Z����O���M���4B3�32���}�	�t��.�A�-螎��Ş�"�V�S����S;͘P8j���+m��6D��e�iWnwJ��V�� ��1XxΎh��>+Z�t���*���_����BH'G��G�����e��\K�Sh$�x/�a_Q4y��ۙ�&P΍�J���"�	s�嗪S�?���Qo7p@���\F�'s������y�=4�	��o��/6���f�L.�w*vH9j�T.$�Q���"�ͭN�k���qT��u^��E:�!���I��5c���+��Τ��GCk������p���w�T\�@%{.�ƎM J��3��'3��2�8H����N�o�t?�r}�pY>��g��6�Pfc�K��&N��V����x?$�&w@�H��������1-�W�0Ҝ�n��7���~A������aꀺq�1G���" c���x�e��)w�	*nW�C��?i���X;�W��m�x�+�i�([)诈:3L�Is&J���3�넮 m�(�dB����h\�]���[F���FJF�_ئ�Q�^��p/�]a�gF�h)�{eb�}ׄm�I���C��7^�������C	����{`8���L����\�����x�G�\뵔�<j9�?���Yru4©J�T����S�"�z�֤�xE�v)��O\ZLԾH���"GS�Ӆ�Y�Յu�U���gٌ�qla-(�>�B3��,2�o(�z��k���;D ���r��<�5��Z��,U��|M3���w){�I��;Pu*��P�e��Z����0���"w�z+��+�!s{���^���5��P�H����c�H��C�=]�b���D.`{�_�V��l˷>Ite�>�լP��#1b��Ԃ4��Ȟ��'� ܄AՀ-�ߦy[�L�*�W��HΡ��z�� �T�/>@^ �'��\4y����,l;�kptdBת�r�Y��/�%��沴�~x�)���i{Ӣ,f�q_� �·��/X��]g�w�Q m�Kj0w�{t���[��d��w� ��V�%)�ʹ�ĀT9(��R����Ck^�q�I�4,�d��6!��D`���&3�&.���D+�`��4<-VH�݅Ud	Y'�F�x⠊��V�Mwۋ�/nU��d�*9/S4��P��D��ͪ\b�U�:��\E����5{P�w1���8��+����q�{&X.����k�E�x����Ik/Kxgb�_=�H�OΖ���,مЦ&=EİM[AR#���О �D��H������<*���\�­޶;�	#�x\����=���-����jnj{`w���nJH)�f&������V:�`
��.��-r鄌�ag��5��]l��?��g��W�i����[9M��x��0����26d�P�ќ��g��.;3��/���-�"Xx�g��6ɇ��y��5>�JMtf@�v��c��_E�o�J�ԊB�hC�Q.7߶���j��Ѝ]����	.H�4ٛ���׊��qS���ۇ#o�H �#�	,�Yk��PeT7w��Ud�Y�k�fp��F�p@�N�j��֧�B� ���1���$��;��@]e!5����-' �{f{Xu/��Rd��!��A� G��_)�._TO��!�95WV���B��:,R�!��%0ކ�q��XU��d��ys}|a����-�k�\_D"��A�I��Uhw��K��@u<�Q�z��"[/��O��۴�2d��9X���ᕑ����(��0:4��{�EL8Q"3���h���%Y+���,��4�H����e��HvӪ+m��0)�v��RΘ^ߨ�'� ���wq��r	3k]�x� �~�f54���ݑ>=4��$�{�1���ai��"�Zʀ#�J��<Ԟ�m{�����Ziƣ}{N#D�k�B�)�1Za:�V�o�\��52/Û٨ɠ����}w��%ظ�mZ���|)���+*�9�s�<V�����57&�K�\	7�]�?Ff��1�w��
`��x�R'F��!g"�ٱʲl����3_�/K4㵢� ����(��b�0�k��u����5O2��oU�<%��nk��t;	�on���	��+��O	!�D;����%�G#�'z�G�ъ��@eX����郝�'���6�c�@4��M��b���,�{j�ĵ�QKE	A�AG*wQX����{l���X
�hRI����К|��eb�x�U�0!i�xb�$O;��1�X0����ĐY��;�~��@N��id�j$�Y�������4���W�M��Cj��u�9�1�[1#ι`��̲�%�:$D߆��U�e�)Yy�tU��R�H��Acz`Ǎ���"������B@���LC[0���U�cj[��A��P5�L�l��&�8��-�.fk��;�tQ's��Rމ�L\���ã39��=���'.�ݸq��oJ��]�aI7��P c��r;�$2��v�. ��^�
���sS����]��
������!����9��h�}4����:=h]�w�~M���;d l�hfS�Q�i�kx�;T�>Ŏ�h���9�z2��U?Uj����`!��p+S.��Ql�=8��b��l��;H�G��o�Չ��(}�`���'vߚ��v�H�Z��R�v�?#d=�Q���y5����%�zWXQy���h���iuHdp�Es*��^�N�n��ϧ������o�r\bZs֎�^P�<|]�+o$���|��za�$�mgC�x�<�q�T����SXw�_2������3��9K'{��*����<
�;�v�|�dpә����k��S�(�Ѯu'8��Lĵ��R85H�;�^�M�^���h1?�V��Sm���-O&����7��b��LzI�y��?�N-��E����2�)^��ȇ��6�maX��0]-�k�ճ�8練{�����{㪒������3� %j�[�Y�ɓ�n��\	��_�������.N�pvw`��l��B�&a��9�q���LAԺ�NĎq����Ӛj%�&����ZE�LI������:�����C"�&o��}^^�R�(��Ea�t��c��rU��ZAt������e^)}��أ9T"l��
j�s 9{r4m҃�+g+��l�k�ѫõ<m�D��׹$�dw,_X�T`��Lh�Fe�����
�òؘ�#O�3}����	/��|�
��.S��M���l' PZڕȭ��!�%��>&����N�9ü%}���+�iHsV; ��Ђ������_�k��
oj~�*�x�:��a�Ğv�9�Ն�չ��iF�����_�v���v�%����^3�c�e1����je�{ ��s.��ȅ��c���=��u��OO���=H�SK��!�!�0.�������g�}](��k�pRB@�a�/sy������17x+Y<N��J\�J� c�bO�N�\���~4j��U��qU㺑L�F�T��e`S?�L\^��Y�,iK�8��E�vɹ@Jԁ�mɛ}[*�Lj�������VN�o�IZ��RkP�4�U�OcH��ZP�
��u�	`M��������� g�^%U��n��>	�X���̼��ǉՀ*�ޱ�Bӵ[�AZtS3�lK�>�0[Ǩ�	��C�G�!��C{o���B�25-����	�r:	�$�O֡wO>���V��O͎�j>s�WJ�.P�>F�?0g9����F�4��Z"�1�c��u7'%��%�ȱD�T~Nӥ���X%��$��� ��W�O��'�:2�q�fGl8=F6�z]ŵy
C��="��{�k*r�l��%�����hw�E��4��ݰ��[���&T0cv)�T>�S�W� ��$c%x

� Gz��:��J�Z|z���c����i�j� 	;V�R�JC���������'�� �E��/ɥ�CK06p���fU��'\��tق���E��j�C=E�^��U0m,��i�<��4�2�[ڋ��(X�����ϭ��xU���h�����(��������m_�|
 `j�t��c~yIc��r4��x w��a���J��q��><�0��Q�6�v��"	�q���V-���ֽ�y��@���i����^u�yf*����T� ���Ȩ+Ձ�_Ĩ�&�uIA�kOKw�g�#����͡�Ə�L��.zC/aC
l������W�OX�
T�p�'���x�Yg��N�/ժ�*I����6\��t�TW\�ץ��y�`6՝�kTUkM�f��Z�'GtIM:�)J�502�t�l=��� ����ȽV� s�,��j3������I�d�%iz�O��ԃ��]jȁB<�t:1�nL�˷��-'92���Mn(�����k��&
V��4E&�T�Y�H�>�E�k�V�.��ޭ�h��s�;��v��7KDڟ�p�\�l��M���D�n]�`�'�:I!2��5��Jd&.�LΊ~��3e����_�}^1��w֋�YJc���h8��I?�Q��"�u�����I�c����u�;�����>0Y�Mgb!|���Dv�.�s�ՠ�E��k�M���?�6o<�G���:pݮ6`	�CU�ށ���t����ç�ݚ��**b��_D�^�ٯ�$�����g�(z������IT��?*5�AGq]���&��Ś�W�Aq�.o���s���w�d�u�4��P��'ё�w�h$B���Џ�}WC'�*t����a��06���U����aj��+�Dq!��yÒ�F��)����ޘ�9��..�����Xq�l�E���+���k��S��c<�5��t��D�/�^��n�m=�+��ؔ����qw�Ɨ�O�n�i��g�v����36K���������+�>��Y�ϣ���{;$nQ�W��|z�(7Ɠ����=x���=$T�/��{�t��kD������\FU	4;���.h�4�3 (������8<'���ɷ\�3�?^|?<k=Ϧorn�=����IQ8�o���vE�C�4���ɛ���aV����Y3]S{ycR��݄�ts(6��C�� ���+{X�4�f_�D{,�6/n�B-'_�&8S<�#5��n��f-=�A�)�E���?�wR*�	��~|6��X4�aZ�4���V�i'�~b���D�cŚ��?:�п�z��"�(u�72��|+ʸՄd­�A�]�8^�hJA9?o@-����@~��7
1��:zl״��C* ��g��Oҕ�m{����c�S�R%B���O�Y
Z�JM/�����Y&�2O�.�my �lv�*��h�!J;�)��������2���`�d�樉�ma���"�vm۬����ų�fsV1b�/��%�=�^�͙��2��S~�]ٔ:h�Q��R@C�Ho-Z'4M_�R�,��Qu��J���<*�
VV;���"߅!��� ���K2� K�`=7�K�aN_�M�����2�z�k3'��n��������thc��I�QW
Ǿ~e��	;�~�FW�5��B��vM��Op��/X��`%?�<EVu*U�v{�\��C=��� |�7Ɲ����v��3O�4�6ƫ�#|zI���@��{.i�����Y�4�����(_��L��n�_+��Ѭ�Wk��e9�ӧ��7/� <۩��%U�����kT�� D�~�Q&8�Z��
�.���D�D�R�
Uט \k��(��Y ����
���7\�/\ �A��\�a�['���>�B�F[�����=\�	p:nJ�3���:s�\̏�8Z$	���_zt�c��a��`Dw�������U
W83q�-4���R|U1��J�51"��k;8[�޳Fi+}�Zn6�zz��\BR>�-�k��h�EL뽔�����wͳe����@�x���h�G��dx�cJ�!�Ş���E��D�
�V�2�pL=Q_(C���h}ʪ�.�M��]�z��Ov��� �Ɛa&�>�?����L!1�Q�ixi�������Q
u.ڕ?���I�����<�D��X�q�(lx��UV�^j+�GX��.��T�R`���.]���{��7� P�/:,�̷�q�~�~/���Қ	�gMw�┼�z7N���l;k��u���y�d�&���%Ѳ��3w��?{Y�-+u��SZ�>b̋�X���D��x�σv]�M���y��xd�� ��gz�y��TS�����
�!^��2ѥY���;B���ֹ�tOi@�6rҽ\�6߉�,�p�?˱=z_G��O����k�'��x���ᘙ��o]b��F%>�z)O�Iد�r���-�$\�I��� ��L`+>pn��EA'�Z�#r�����k3�����n��>:��������� ���ނQ��QFݷ��h��E�JG���� =[R���@j��9kl��0���6v#G_uk �>���Uɯ)�n�)&���7���;�C�e�X�\qG��N��ʤ*$����E5<���v�1�Z��y�fUy��V����{�#F>����*!5׈�6@B} T5�n����ȥ]&Y���^�f������OJ$qD1��V�2LaY̦,�x	�OV��"xۆ14�����Y�.����c�� �v��Ω����16��y.Wơއq�H��׋\) ��+��J9
� ��w�)� )g���3�p$�z�2��U�x0s2�ISh�5)n�~w�h�Ӌ.k�V��t�f	#g�dܯâ����'�di�3�b����i��"�����j�G�Y¼�p}�
ܧ�e�F��f���B�A�q��~ ���th�=����3Ө��fG'��׊Z���Әrg3lsI,ёE{�0�I�����oy7� V�iN(�j$t~�|L�&�_^���S���alwYy�=iBj�&��9�b�ț�5�?/a�ks��Yꦓ�G���!����jjv�����}4�"j�N�JwI�N���r�ѯύ`�����=A&��pn1Ig�EG:i ��T��d����1���W��4.���qŰ700=+\��ʶǭ�&�<��QQYl1#���P�X��`T����'�(� p��j��m\}c0�g*���u3TT)���'DȄ�=)XT&����;~VX�{� �ڧK&�k�03�y�on��|�b���utV܄A�¿� ��JfKZ��P��n����vf8�����Xf��M�Όfe��m� 8c�	��Rkl��9gMO�ܓI��3��?J�ۯ�:P���T��D����n�����8�R�s_�Ѧ�)4`u���)�Fu��X>�5�!���#�ϰ^n�['>}R	��!�w�fU�:�E'�NM�Y�8y9;����)�Aܴ�?���@����RBM(/���.��9p71�2�Qگp��7B��b+g�%+��������������\�4������;w���̳�#[�6���
O�Q=Ϻ�]v'��JF|%�Z3:��������P�Z�2ܬ��|�nI��VT�2>�.F�L�T=Fth��;S�$���0�
���g��9��H^��J� 8P���k�����Z�L ���U��eoZ��,���{��t&�ѕ!�דPC
��NH���m&��ȱC�1֯�n����].B��+��3���-x}��*�e� ����+������,90-7{a�7a��{dw���8�IfF�������/N��� w���8�"R$iU���H8U�5�r������ٞL�<-?�*k��T迣$G��#�-q�Ң0�
̩Y?����B+�#�2����,F��ʨVUr?u
V��EO�cF��X9S|S�g{�$RK�X�0>�~sM�_�l)���G��n�}���T�i��s�4�O���l��b��X�Bl.�XzO�O�^<�����3B�<�T���Ls��!ա�j��.������KV�QG �疫�(;CS�3'���<o���C/B�kK�R��vwL?~.�ƍ ���T��%�Q�K�xyX�'\��=;*�����b��~�%�\��Ѡ����?���+�L-?�X��Le��q����j7���������2��_6rG�`>:%A�W�WKÑ��P�#,�S �(�/�����g=I��C�e!��C�U�L95��ډb-)�+��D��`/}{L �Ɣ���Yz����+(lL����L�i����d�y}ߨs������Ʊ����,����e�; P�1�(0�����5����W�u�t�NM�(�[�>P%���J��y�&?����88a��F*�Hl�y��E:~��&�$����;L���ĂQn+x	�.��Rr�mz�E��?ģ���%q�~�"4�~�Y~7xfDd�J�����Y��J/l
����jh���Q;�lR/z�-���f�E�m�x�����ni-��6+�sV��j^iM���9��ʐzM�O�܄��"F�f.i��[�!������L���O[򾹿0ޚ"��H-�3��/C���d���}�y�<��X�-��PDhcUC^��|#� �>S�m�(:�+�� �TRHDx���rp�:Fu *'��Y�4M�b'���Q��V��I�6�B��&	��|�.^��E����x�Tz8RU��3Μ8�2���ߔ�x��_�W��Ƣ����utj�H��̰�>�y����P*H|~��Y���Q�(�(V��jR
��QJ�yv�4�� W��`�J�Y�n���pX�{s�ˬ+j�-�� l-N{�r�l�>���y{o
���ɋoc
���f ^�����1���I�%R������(L�N�pŀ�0�!#6 ��vc����X��c���.A?OS������O���ʳ�x���$0�b'h`|Т����G;Wo��K�SiC���"&�TV��r�7�i`�'�l0�]*.�WB��DA:�\�/�/�"�������&PF�@��=٩�(�N�@w�*��:��ᜢ��K�Δ����0|�/�%�,��u�a��j��ۨ�C��7��$vw�o'b��J0�T*��?|���ƌ��|^A�2���j�".yf�CN�6��!j�E0����E�_A���5�\��⸩�@�j��%=�k�n��"���q[hs�k����~wN�m1w!��|�?S�xȕ,t����
T�\:^���^��:2�$�N�k.˜����b+5��!p�t���Mc4*dQj��͐o|�~�(" �9�eC[��m�gg,�SQqOre�Y��D���_��V��o�\�Sy{����2e_�B���KRt���N@�?���A�j����,7�miJ�(�)� 33+]�;�V�^���C?lj΀#O/�(B:����y�gt(9d��7���o"@Emk$�v"]��\�ƪ>hؾ �ў/�Í<�<XI-	t��޸�<�7s�IYvD� ���EȤ1�Ya�}"!'e���M�<�?y0/�B�������պ?��7m5�qWH�_Z*�CqĂ͠q����ʶ�	�Wc�u������Cmc��W���J8;`8�ȋC��s���	��t���g��L�]����L�Q#+���3Ϟ[� ��Nb!�,�J�����`�v��~�4�(SHM��%�3u�h�!r����)`�xo��E��~��8�H��x&$�~ 9#�@2��t��_vGfo��V�ĸ2&��F��8��zP#R(��#�6R]S*�{��up�8�*V=�'E%�>�؜�'�x�4�>�E�oF#CßX���k�vS w���б��k���ܪC�$`#_�2k-m��)�Yh���u��=�5���T�M4�¿�V��#��{,�P��rh�J;��Ơ�,��3B�2�vW�˺��KP��q.�����.GZ��>Q����
ⰊD�M��"����/M��W֓�F$z����7>�n�j7�	Z����r[�g�\;п9?�-�!NѬ�D�8q
0�gv*[�ӽlA��q5x���wx�s4�a�Ps`�Õ�������w�+�|�O�;c�?��Z�zH�@Wi�b����O?,�{�Y���/F�)~�O��UX|���^L��Ns���R�?�.�@�ف[��=l���E�]�:i9�2B���1w�G�y�}�����:e����ik� 3�޲Y��K(H�>�Wlz�Co�u�%�qa]�헎XjD�����c\m$L�l���ڑ%�7ڨ��wbz ��� ��.�9��eA֎㉈��Xh l�A�k ��Jqѓ-S?TWˢ+L�ߓbw�;B�Z�m�g�r��&g<�n�0yX���Oq̤��jqz4_�ee�S@ڡ������["@ ;*�]T��BAU�PT��K�{�ʢ���1���!�2Ѥ�/3����1N2Z喸>�kf#�=.�]ȷ%f���������]��r�i�n��4�EU8�~�Ejh��uSC��`�5Q`X]�؊�,z���8mwv�@
������d��&�o��u E����8�M#��3���lQ����K���*�yy�ѕ
�������
�he�oxS�ρ'G�� ��"���1��?��j 쏁��N8l&�:�������5)Ӱ���L!�H�gv'�\G�2�y�7�n���f�l�"#���~t+^ `�D,.�K�,���3Ah��l��X����M�t}�1�3M��G��V�%XvA,_#<��}AG�b�ۮe��Q&�_�]�<
���!��T%k�>wS�N�ƜD��-4�ř�}r��R3�G�1�w�څ[��;�E�A�L�w�뵃�y�(؆�Z��z�����iU͋�B��(���&���/�F�	��I�1��,�b�i{_0�e�1��hH�v#~�b��.�����:@�s���j�A�&~{��𿄚o'�B�8�XY��e8�V�QB�2���
o�/a5�"(�Z������1IW������ώ�]��cE��wfG�������|�5Н�H�=I\�����4�mk�VI����`�Z}��K���H��"��.�nk�!�����#5k���
�ɼP��XK�����08gV�)��N�+bSC�F�`����v��UY݉i��� ]����y_Ŭ���{�]k���Ou DcQ�x\e�TZ��zRE$pI�*R�Ȃ)4ꇘ)3gق�t{]4H�k���L�C���"��c� ���ED��e�L���#4j;��q�J���v҇�S�ͬ�ç����h���̶�e�������io���.�~�����r�|68ւ�vО�lѻ5d��NUᮣ[�z�m�$t$m�~[Xt����5#)OGG@ؐo�(����7"b[hwOe`��7�mp3a�}z:.a���@�>;�`8���u��<]}�~��ǖ���a��O(X�A����i+����
�CF�a�$��Ѷ�vL�\�ț]f=?�%Sq�of��K�z��R�H�8��w>���Fk����j��	�������Ĝ����X�@ͨp�i�<�����������g���U1U�cBZ�ъr4���s(a�sP�I&��V����E_�Μ�2�����F,mLY��'i �����~���K��~{�Ei��z���k�K|���*��3�J�����c���)�j��ԯI9��eb�G?I?q!n7jO�qy5�[�{�3��`$B�m�_҉�e�;�����7�80Yj�׈AČ 7ա��ѹ�)e�=�.�h�e%zI#��m�U5��Ɵ����9�$�[��QZ�)���ٹ�r��-Յ�^ �
̃�)����H�j�a�l�(85\V��g�tJ�wR��˾�}Xq6�d" ���䷷rX�`_2��?�+;)^5��L'$	 ��/,���G��>���	�1��!BꣷKP�-��I�[_�lG���·����{�>uVKCnu�7&����#�Zy�{��-�':ұ]�A�;��h�kJ`���q9�(�㥢-5�= 	ꌩI]�P*5�e�w��]�>�1��	��yC���S����ݺAY�EK�d��c�ԭ���\O���WX��#���k�:y��N2�kP�a��,BF�\}�ƈ��'{�C��<��y��UQ�j2����r�>bL�������v��
얐��i�D�;��%n�M'��yX��YB�9��o�s�-~�0��8����aI�|��	�|��a�߼\��s�uQ)�f�Z�ls�56�5��cXgh	���F�$�	G~�̂��د߃�XC��,3B��+��-���J��g.�4IX0ʮt�o���^�eI��Gc�۩�z n�ݱ�%�:@�����Q�W�·�z-�5�Ec�@�����Hq���4A���j��n�G	����}�x��L*ز�p�8�Iч��&uB��b�:�
��P�WJ���2������k����`ӊ�tڬ"�ef'��C��p��:dG�'��$1�0��^`B ����!�NA׹��SA��ɘ̽�I�Q��a1�NmY�4�#60�Z�E�U"<ܶ�N��n#-rת_r����I�ׯ6<H�ö�Z��l*�ڋ���Vѩ�b�{:N��5��R�"gX�-�߭D�#t�� ���eRʿ`��<u7_�]e"-�7=PsúA�8����g,�H��1�����c�xbO�ġ`��T�F�9@��x���?H�\.�x��ƿ�{
K��z��+�x��q� |��v�jyA�=��瓘������4r#bʤ���3�ph�Shu�P_Y{�U?��N=C�n�%Zl�|�x����Y��vEV��1$;:�ў4�V\0
0�w�X��h{�Zށ#妆���\�W��I[9��4���5�V���_R\&�Y��K.��)�i���L8exܤx�fE��0���!� ��Ŭa�M��G�ťy��:t��ݼ�/qԝ�\�Hk4O�U�ܿ�k
�S6�L����R��W�VG�%� ��'7T^�;	=�`��x�W�ocE�#1�쐹�d4Eӛ��m�fm��ؾ��0�6f"<��n����-���g�_#�k�Ѿ�6�i�]������04�2� z 7d��Oeu�~��B;��N?�LO��4��Y�K˽��?7�8�Ia۹�⬌Ţq�>~�;2�-p��5C��5S�۫��򺃤e$��4�P>t�U����8M��)����Qxu��1�%ޫo*ZV�9�B�E�#��b {N�9�l5��ϋ?��H��ǟ��S���n=�ѣ���3��ך���a̀ԭ<�N'����0�H�ze��ު��/���������D� :�4ZN�S�.3�,h=Ou.W�Ul|ɟTĎ����uh���׭n� ��wvr�n�q��Q��4�u��8	<q�6�`N���Pn}`�(z�g_ׁ&J{�S�;UQQҨsc�w���s�#!bj�.%�L|�AǵM�BI��1q� 6~C'�����Ea��?Ĉ\KހO�� �i�b|���/(��Z�
�iL�֓�����_^F�ֶ�뱼�6��L���>?���z2|+�³�D]pш���w����Ob�F���
\p�/�R��U�rp�Y�g����0�X h�{X��,#!����u\I&�`�`33y 3���xj%�.7�}����j^ܩ��TJ�eM���"�hp+资�ƶ2�[�"cXg��t���������
L�k)��xfd-$�=��ϒ��н�D���Vj#��c��zZ���T��5�b��.����P<�|YI�9���7k�h��V9�
����cF�hqġ����bPɘ8�v�����Gâɇ� ~�x���2�|����@���P��6�Ћ檭�H+IusǤc�*��V�'늪�.F^u7!�3.>�tj!�p���r�ؾ�`����d���^t?<����m<��U�N�Å���{nc�;�U��!U���0���岵3�=�$	�&2�@F�w�)���Ry����ʏ0)�cV:�X�'�����JP���#Mu@��x�F|���?M2��VN~�����x4�)74�9��7�!���H٧�]xH)�e��s��<G�������鱡˂sI���@�Rb_��3"�\G��~%#j&�,88�zXc�8��[׬�uS?�-t.(R=?QG���M�Z'd�����o��J���_�&J���Rwתf���[�b�)	M��'О���0���^��E��荑;����
+�q�F�T�u^�Uɶ�e*�<�.�[��	��l�?6w�̣���/��o$'�S�Z�}�=A��֞T������Ѳ��>h�6[�����R��ܮ�ͽ���utoN��[���I��M�5��.�PF-PE]k�h�1��HQ�ة1]��(G�4D��<R,d���0�v�����䗵����;��ߐ�����o7(���0&�(�-2Y�TB� XBz���w*���<!�����F0qb���M��� tB����xb�ﺌ
/M4��w4PU��lY�0�'�{�d�*�[o��Չ�J��z ������0}Ƞx�lE��Y�����S|�S�+�]�-!����J����L����؆��b�pF���IJ�K<��q��tQ9L/Q�*�=$��^%RN�f���x��
���
X��u�P04)���[K,��J�Ye��(��	]��͌�Q�M�|��Ey�u4�\$�{�WUhSh�v�n�Yo��z��z���̦#H�F���uD �ɳ��l�'�Eu=AUH0�8#e�<�L'q-�E@��� ����W��e�I/�*�Ւ�`̢���W�b��UL���%���~. O#'��iJ���}��C�=�zJ��~��m�,@��ul �����M�N	���j�N�Ӿ����7W��)9A��w-T�߂����X����g��r";Z{/⃹�e���p��}CZлY�[�<�I�˧�F�#*6��z�i�s)��Q�n���iْ�������/S|�/٨W�N�j��zsQ;��KV��n��n�\�2���I���S�]�H�ꈷ%��Q��Ja���cta�W�6Bj�����IcaM�aW`��m;3%��t��1XO��%1C;�
���❱�U��_�[�����Cɞ�VՑ��j�>�)&�VqF9��L j��Q�$LB^¶�5fD��I� ����*s��t�є��q�f���R5��
��HΆH�	F}|%gE���"Ḷ`�v}��!��?:��}Mm������yr�0���L�W��n��4�������-N���v�c+��������`���f�v��:6-n����?k~0��d��49���Be��J��-�: ���*+(EfJ�8jDj2t~&�ˋ�$;Yeq����ă6���W
1N�)18��/�q��R֓p!���AS�̢��ײM�6���JW��0���ǈ8&*;е��U_z�,\�����Ñm�p|����;Ok�2�9%��^5���C�IMI�%����@ ��.dWȋh��V��JBy�RK"qjq� F��:�~#����5zi1ᤛ^�ً�x�UK�?4q�߱�25�5�7�^!3:c���M�z� ҸP5	�9��;Xz�����:i	���u
��^J���u8�/�`듛�I��X�����~�i�%�r�6����З>:��*.��2��?�"���p��(/��;`vR]��'�r�*���A�P�;'�mIr�B��6��4�N�� ��I��PK|݌w���
^<�R�+��3ӗ�Gz��"��2X�fq�}�\�q���D����	�L�S��H~k�7J��-�+�7u0t��m�
�:�!ೀ��Lki�.�'�P'��^�ز֗�j�<�q���+>毄G��qQ  '��T�@���G|'�o
����n���1�����6�WI�����n��5��ؠȭ��Q�r�����y(g�g�����c7�um��A♌�2a����{:jQ����9^��v=8reB �)�Im���Z��>j�x��9�$�t;A�+�;$D�[��T����S3��'����qm��
.Hy!���e���qX�؁g)���v��33����q6��#��)�=c�k)���(�CdP��@H-W����y$D��@�����mM�x-)�0�a�]�ϳf���I��i��y��E���2Am7L0��%`�)���HK��r\n�bhr}��ţ6Z��{D▏��|F����V>��(��X�|�R������hE�x��pGgي#��,Rq,�S����=��^����ȂR喺�h�h�/}�8{�&���l���8�2���p��̽ܪ�f2/�;v�V_ij�B���z������[�C��/�������x�,������zDh?7��&eM�i���\��'#H
��@Ț�L��4��`�|�7���W���5���]��2�a��Yެ���',���Ec�溑�l�AgA�^ �e�Q��K�ґy��>��
l���1f���9�U�ʱ�l^Ie�"V��&Gv�+�
\��J���^w���
�	n�;b�;:�3�V��rTؖ�����m�؇h������W
��@ �N�>˔[i`�	����E�6��CY)U�I�������S���'4��R�C���Z%wŧL���L��U�B���e�B+ ��cOqU������~r��)�~q]K�iU_I:�4yDR��!:s�Ή7�%a� >�����9���)\��V�w��R� �\Э'�v���I,f�Z![�B��z��%k�c�5A���B�SRZ<���$�TkI� g�:�������6����_
���[O�s];	 ei�M�K��?��w[|�L�/��a���/ݹ}׏�!��n�*g}~i��)p��d0z�z��i�à>��$\C��I�&�$�yxR��Cb�9A�|ژ��w%v�'��x�ِ�VU��" $�1�+�ߊ�1&��h��e�A����Ό�*Р��c�~�!!l��5F^��s���y��o� ͐U�zxVF��
������w���׽F�ι��q�'��~� Hɢ���T�X�H39Ц7h�֜�/���v����X�q�8�)N'��N]t2�E>������2���Y�D!��RTA�)���࠸�iG���91�������i��j�<���U����K)�l̀�b_�O&�d���}���o����������j����\i�S����z@���m�Vd)����'����\3M��´	盶>n���.���{i��ECF>�r&zY��N�����2�#��m�s������P$�ז�^��wɌ4B���-lY�lRL|�����M��`���ɨ0�}���b�{?�̢`�1\k5�����P@R^���~Fa8����1yQ?bl4D�2�BK/r�5��2�C�ڽ:��Mq�W�>Z��m�ea-3���S]��k�Dh��/> 3F{y]�T��9DD����_�Izs"t���4�i�s@��69H��%�����	P����o�-��Q,�q���F�hh5�w��٥���5A��D0����U���6�]��l��������ϔ�2x�m�U��ޭ'���O�t����L��`ZQ�F��&���X�n��%22�x��"Mԉ-M��~�	�a�0�~���2����������i��J�ժH	�Y���$B�u@��e^e����x:�-U�gbj!٪��#�9�;�8l��Ĕ��KlJ@�x�Vx���tY���T���a܏�њ�D���8��4Z�e�d�[y��@��*�=wY��A3��J[�YΦe`�&$�I;�B���cV�'�r/v KǙ�dɻ��l�P]傫�q1���@�^#�:է8�iy$֨ӭߨ����NfXy��~گ�:������Y�U�u8��u�~�����lƊ�����&]�0jZ��B���e�4����vPw?UW���6Ma��'x�5q��:��;Q6H�Z���C��A|���f,��[x:Ѳ��(H"��1]>�)�l�C�{m�E-�d�ڗ�x�)��G�%~b�,X�7�N����`����:�oa{zq[����QR��ק�Ɵ�A�[�$�{,������k��i��[^,���}��oe��b�W7,�)�H��Y;�9ޕ�����cWg�uʵ�s'7�P�Fh,�M�U�ա�c�E�<8��{-g�)J�������p��;�����7F����y#+��r�p��1T������hmYCF�o�\�����K��U�������S.qҝJS.�6%�e���̘�b��&Qe��S�נ�
bn�E*=?F����z@?m���GD�q���C��z�B�����:~�^���}�n�7:`���ӊ�[C�(�E%���?5Ϋ!��Y�0�:=�7[+������.���\ylg��^�'�oV^���9h9�;��*4�R��Q#�cJI����
�l/K�>�"��i7���Yc$���S8�W�q)�I�=1�Y���'n���Lan����O�#�  l ��Ȑ��?�ܤ=�gl�s+�߄�	�K�N�۠��Q��ԗD��\��FL<Pk�1���Ȼƞ���,U���l��_��������+��$��>�>u��x����W\h�m�����롿���~L�F��Ǭs$���N]�����g��I!i��`l{\�8|���:ހY�^�8Pt���z��H+�	��A~}'�-��hJ�q0��j6W��"��;��{߈��tI�"7��Hh��?�f�oW/���X��6aF��#�4B�	�����O�%�"l�R�Fd�ӊ�xA 1��/V�kV;:����4=wX�j���.�$i��̆tB����u�]а�ö��ͅ�YpydQ�
(՜HE�:��o�iP�{��yK#�E[����S��M��߂�����<jd씶�T�]�E�0]�ƶ��8�|�W�3���o�|cQ�`Lm�]YĀJ��6���wk.���h��uM=��b��A�*s&n���Ϩ�N�@p�yӉ���m!�c����ƺj	���O@�\DW���t�NR�Q�S]�o�����i~C�[ ЍB�.�'�o��:G[Oo��`#�es��'�H#���j�{?�oТ����שl�h���A���U��eꚣ��V��&�A~Sd�E�4�S��R[@��� ��c�UP��NMEw�1�CM5HOG!��-�t��!�]�uzު]�N��
��<�ގ�2�=ғ��f�`=�J�I���9�[O��t�%`��X�p(�{��(b)�)Mw���u�	���k1_�H;A�
;�I2p��UoWSz2Y�C��$-�����*	�Ϡу��l��s�e:ëg+�4��C�����h���d&ߜvx����Ə��_	ݽ���%�BbR����@n��*���a���*�tEs�Sk�������}�c߯�j���'5x÷�����d�,�m'�9��n�{5%����i�"�Z�:_��+����Ti�`�v�aU_iDP�'��GB�;�2{E�	����Kpq�{���m&�� �]�B��\E}�9n>�kT��\yn�릾o�UBY��}�z^i�Z?e�>1r�d�{1G������X���ї����EQ���˜�fgp��:<;���>�w��r�#�T�����nzA?�|'�xɲ6C����Pu�%{zF�}~!ˑ��5CW�H�b63�,@��΄�[�.���k�3�k�8�a<���?�~��x�|M�A+	�2'�A��>�j��D��u�ճa��5ֽ�LB��w4H��|d�<̓����1YL�^aZ�	�:�S��ֈk����p;C������x;}K@%��= �b*툑��V����b���~�%�W��f^M�ƛ�u�(�W����W)�[��)�ĺ���o��-�Ka��q�xۅΨ�N���i�T��ѣ��b6is��~"`5F`��Bx�4�+sai6k~���Ŏ:���g�[ěk��_d�/<
+��D�'���������-��)���;�M:�kbЫ��ކ0t]V�U����i������=_e�Kvxu�,����w&Y�n���HY����˺�-��l�J����|�dx�{�o� 6���t	�_%�[�<��ޏ�K�(��A8�����6"�<�o����J;�V��G���`�o�mBg�S��{�55�D=v-X�ttwLhf��I\��nc]$� �۵`Q2BnfS�o�����p���~�N �0��Dm�q�u���K��Л��\FĚ��'�k��_�G���,i��@���~���x�)E�ϵO@�] 3�@����%`,�1|�&�[D9��|<]�zY�m�6+J$X�u�d�W��\
>U�s,=y�V�Q�Y�(��+*%=�����Ͷe�O�Mdf@E\��3��D��,��ʕq�ih��D6Ѷ1�2�/���x�+b���F [ب�윇UJLs�rE���^G+3d�uw�hVor�ѣ!�,r��>����z���u�y��^jtW�ʛ��H��Y�XT�7ŏ�C*�Ԑ��k|G������vk�OX�-U��;eR̨l�� P�'?��t��O�&����0�E�C�S47}�m�<&Ϡ�tjyLN��<T���LuCo�rF%z>t˰4s{~�~�;b3�9D�j=NW��V��6�:SU���"�G��Uv����{MZ4���t?�:h��?�q�4��tTB@zCt��5�״7@���pwձm<�_�u�LeH� ��&<*mrў0�a��D>��.�.ռ������j,'7K'jC�bLh�6uT�����O*1��'Fů�U�}�����^��1�5zOIkhAM,i���P5'q��ʹE�Ri��A?R��\	C���h7���#��Vh��Y�'A�Q��-�8���	�ޓ�Hrfe�6I�J���9�h~"���.�v�*GK��2	���`wD;".����ւ_��G �j(_�m�Vuj��O_���Z�%p.ab}+e���Ä�2��Ơ�������y�NM�v0�,�w�>o�ԟ	|���dׄ�(ۃ=��5��S�uZ3.g{	n��d�*#�
��å��~EF��?G�7�3���o��(��QMG|*�|�u��z�ͼ�����%�S>�O�D6żKl767��s���z�7v�	%�ƚ.;q$8Z>N�
Gd�ٮ�����&k�hؒČB����t�?��>Υ�������>L�����D0Uڄ����[�Ǖ��7�z0�~*�5瑰�?�|��O���C׾j#榎'���%K"p��� GpXj��I�Hx)}���ߊC�Lj�u��볿�f'?�>$^��"��X]�v�\� 
S�Н�=dt���K�I�ftiW�z���UN<[れnjD�c��
p����Vó�?�/�_b!KT[vE�E���>��\6�� ���LX�8����� P����sZ��u7D�Ȭ�!��J���RDq�����B1��qXI�a����Ab��Ζ'�XD1�!g�f�z٤�%]:�Ȣj�OHr�f6qR;6���r�H�:��˥}]D,Ηq�7JY]L�},f�1��"�;wė�s�Fn>�KΞaY�Yf(D���uJ"�w�T� �¯$�3���kP���=H�}�'�����x;12k '����K�IΜ�H��+��A����OQ��c���%_@;�7E��{mD�T�Ƈ$(�>�ǝ����u�ש��x�)""16��6?��E��T6x�~}�~�<��e��X��W�4'b�ă �C�p	��$P"�������O��\�ɳ��;��W �yÀ�	g���l�"�D7��y�:w�ye���ko���ZU�[��q��aژ�%�O���iD���`��?d��ñC��յ�����Z��@��7,q�	���$��ނ�yۺ l�XxD�=S�"+�9�X��l�x�4ɰ��ǽ͐�zИ�1��QYڏۤ(��}��W`�?[��ݼ��a�7�?�h�����ρGP��h�-��4>�+��&$b�Eg5�����˥�JM����b�}��5��N?�9v��22�����A��A�W����1-�XM��Y�$@x�t>>nX��x�
���3:�P��졻�!��io���$."s?�v��}	���y�NA<���>��^�=�W�k�er�ì��� �t�g�ǖ�͝t��� Z`��~�2��M�<��݋���;�B/GD�1��_�\�a�n>tF����`��J�ޫ�[X��M����U�I<��el�X�~O5�,���@*�p�y��;��{|�_>{��w�Z�,��e���RL`�e��6�Z���owI&�#�&���0�.X�f��:ѱ��/q�+��!n	:?��-��I��X��W��?3%��B��X�E:*�9n.;N`�D���H3��#��t���i�.z�}\b�7�O)
˟�Hq߉��!��_9G�$*4�l��R����������Da��;���Y`\��O�:,��pX��L5�?��D��~F�)�p9�vSF#Q�a3H���S��ݽo)G����45@�1&ɸ�Qfe
��6$��-\˰�J����J�TMb���wE�yr���
W��� �� �~t^ێ��h�_	�G2A�1e�i!ĿY����tQ�:B��OL�>��$�*����ؖ��k�v5h޸�����Zd
g���TP�]��%��qL�Y}i�6B.�fi[����v�4��/���K�:ߌ�����}�Y�ςPO�wcաÀ�O- IɞP���b�
����YGw�ye�A�bĮ�	����Ui~�9��>	t=jWS$1��0��O?�o;�����T��z��G~cI��:o��7�e��Mz��n��#�R�Q /aM7�JO�`?���{���`��NL8�	"ʑ�4�Y_� ��,�6�Ω�g�\
_��+؊dS&������2X�B"��Y�뺎{`�U�袭eB�©B�dc4��3�9�;`% ��m�J��y�����-�mT�\Q��kQ���h~��X�h]}���*�(��6�$�'��G��隩Κ�&m.�E<��tm3�K���?��J�P��bG��H8�; ������Hל�HF��܌���>dO��M^�+�>E.^[�¦��%V���H?xn��_�[ �_^�r#0m_
py��*8�w�B��2R=%Ï�Wh۲׮��]��G>�;����O1��s~�ɬDE��Iy/�L5�@ �y��''�^�ؼ���(V��(`���N�����;�NA	\�<˚ �9��� �d�QΖ��Kh�>��aN?o�7��(�p�s+����U��6�r�F��S�ڷʺ�H��OY�'�Is0]}�����i�X�Ʌ�P����2��q#�7�w#ҵ
��8^��!R5Z�j,�a9�Z��ް`�F��ۈ���.�ٖ�$Y	��آN������5�58
�T����������1��>���U��`�0]߾���cر���k����ņ�$%ݴ`�$��t��<��C��l�_�IAz�o[_�	�����s���`�8 Ԋ	�a�c��}����)m�_y~j/��t=x��W�+�ᆣ�h_�ɦ#�Y7��_g�w�����sM�.�d��A�@r(�ŕ &h0�<�R�?������J�r��m׍I3ŌfoG�,Н̮���M�6L�X���g�N]�yLvqv����8�R�z��ͺJQ|Yp���'�B��l�:PrB�QZ�
ԃ��L�m�����\�ܢ��Q?+���I�'�������Gd����6�N�7�5�=k��9��v'A��ҒY"�Ʀ�z��Z>�f�Þ�چ�MW����9�w�['�h�-�.��$�C��;6ܞ�/�J��М��8���0k�s��!1�G^9+�j���`����)�����q�O_�]��I���N�$)�͇���V��l"B�Ċ";���ƛ�r`^����b#O��K�|)lhN�����x�N �\q�����6�IT,b4Ϳ[�IP)��zb�k��&C��²��w��m�p����]�(}�l�nQYd�P����ny�'0��k�N���G&��-�������H�Vb�0ǯ߷�2�Uo�M_T���3���)x��;��8�rԅ\���-b���'�u�����6�x���.�Ds{.'G����0!���c	UMX��Ép�n��Z~*��V!(�y�N�)x`�&��#�' �&�����S�� e�rPG�mUuz&謡&�4}��]��r*C+��OTR�D�zC�~z�d�_��,Le�-B.��f2�;�)��*��N�h��x��G4��(vh3����Irg��!���Lc[�"���7��;����H�����U.������'�ѷ�֞�p��}et�;��p�f��?�{�Xeq���;�=B�R\�oʀ��H��0��\u�%�����H3���3(vIh'RA����b*#ȕF�u棉�$�e��8�w��=p�!��4����Ƀ��x�5E����q��_��a1�N��lPo�E���6�������������u�+%?x�o��)�,�m"�o���%�i�
��'��-P�w���-mt��%��@p�*�81��5ƚ�5uZ6�b@_l`/ �
�i���1Su�2083�Uܵ�� iZ��Z�>G? lm��*��6M��w���\O��ǆ��vD�Vk��čz��hч��q�?c�Jr�2���HLL���C��'�/;f"�[4��{��虋Eh
������'L���."J�bT2�s]k[���&j�LQk��D3�����b�L��d�a-Z.�CS:`�Ѱ���o�_��1�MSFw��I��"߉K��zE⼲��Πq�\ꃠjz�s�"����H��Z�v�Px�v\���XѵP��L��1:؉�*r��:ALb
2>�A:����]qC�b����MA���	�	y��
�@��fWEUF�!�OI���E���Y��:;���S�t��{���Nw��PYn;ں��V���7Jp�����OU�|�M�e�Ez��O�Ӿ�����=-*�éu���Ώ����N�7������:˪-5�_ YӜ�1��Q�z�~&7ހ�A=�o ����,���m�6�P���$E��d'BU����>�4�.��]/V/"d�j����0�T;Ծ�A;���ա��{����@mX_738	���Hg�M��'qFxY�5�?�&-?}2c�f!&(��|���C9�u
�X�M�	s�z=����b�B�x@yO5�#JK���U�(�(�K�����bs�dE�!I���`���dW��8��8�D�~t�F[���Ϭ�+#����r�'�\j޽m�_Ey&F��p`c)(��y�HУ6�-
8��P� �����6�eD�D�,{7:�G�q%a.|+����~���>�QF9�����`�܌R����������j5+��ٝ�e�f-}�p��L%�κқ=��V:�����BX72V\}l�����L�O�s�!pn����њ���PI��xb�@�4+�ȟʕ<��7��ԳB}[05��`_��[��ݣ���.����U����pp�	O��f�W����GW�AP�G��vO�d/��u�RioNirå�P����TkG�"�p~�f�W��nP�}�1C�g`��6�xK���+��L�(,�iN�߅�m��Ǭ7��9����b�$�;O���r���9�ܾM(Z�8e�Mg6.9�&N�3�+y���, �k�Z����D=��YB���@��h���yD�'����z����K,�,/p�K7]㏡R\J�h�c�XԱ��~���|�P����7溆��f] XQ�]�(N��)�m�;֍�|����~5j��־��a}�Js����hD�<t���q�m��̓���@C���s��i��@�K���9V
+;
�0T�+.Ę�4��	v���z���Q^��d'~���{����hAI�|�uKL�I���ʸ��8�A�X{�N��Ι'��{��H0�*�qW͟>�7��*���ـz`dW��<�7(��J
�|��J�h:��C���������7��7k`����dEd�>Wd㛣��{��v?Q`��M�4~�E�E�K�B}_��<�AΛGw�Q��
z����My�O��͖��V��X���e W��Ch2R�/�ī��	;�>�ȁ\5ESz�Nj]��8Hm��3d����[N�r�{�E!x?�3��N��`�[T��i��RB�"� ���3D��w��� �G��*;G5�����7�J4���������T"udș����̋��kH��,F�*���`���!ř�R�}�Xu6�2�grrB�UϙY��ݠ-�3�aq	�W��N���&Y{_�nG����k��\����qʪp�-A��D����^���u��[���y�o�l/G�rj��������WJ
W�e��[���æ��W��*�okS������^"��1�R�.ￏ�^�}JaF�Q��@�D�$��	1�0�s~�d�N��/�Zff����_�G����Ϟ��f���^jd���׳�ţ�H,���� ��G��|�:)��8�N��� ���2��fF;�*�?��d�� yuk4�+�9�T�@��.���6l/��S.��6��I��0��GD�Y��������X�`�Ҟ�E���2�!�X�\�HO�')ޚٍ��b�=��Y�V\��;��.�7{+�e��:���*$�5�1��/B
Ůw1/^J:�Sɺ��0�!�mϦ"�o`��]pA�����g�"���h��h��&��U�ݤ�����,���!�幆]�Z�����h��σ�7�0n��׿�CEJ�GC:�0��`鞆*�]��(�,�Tm��3D�`�q;�@,#y|�)�����_��`_T^'�,�<i�h��yrV�����,y�
��=�hB�eGgj	��z���}x�e��:���s��૰����C��!�k�e�D�M��RB��B"6�����27�J���&h�+��!KN9�������HÍ�;jՊJ�j.4����\[
TOߨ0��Ub�1nD��9�ր��^i�T!��P�goa��[���;� �Q�cҚ�X�§;g�����Q.��>��tB��EJO��ǰ���\�+٤�0����ƥ�+�hl%2J��(��2dg��:tp���b`��`����;
H�yk*��]6��`|�x[�L&Y/*Xӊ�p~,W�/��=�����LW��ST�����EW���!p�R���~82h]Y��9�f>Ϩ� T�v ���y��Q(��F3��4�;�_W��(�Aj3	�=��q#�~�{U�G��Q����(�ksE�Cv*~�����ѡ����,-uB�M��:"u�#�K��ZkE����Bve�*���[n�3b1֒HavM��ʪ>����^��މ�V�Ӻ��_�.Wc�ަ^�|ʝ���p/�ux�J	=b���YJ�C����D"���+�.P/�~^�G��ki�u)P,�,��y�����6�F>���:Ո�!�hJ�O��6q[�F7�'�F�R�ֳ���V5�(Gw�Zգ*��}��e� /p��Q��f�6 *��n�[��Qf1h[$y����Rc̣B����s�g}D͓y�|�=��U�/O�H �/;�KǾ"3어���ѡ�y������>sm}��a��:���b��͟-�]�#���=����Cpߺ���>�!c�)��!��6�8}��0�\�G��.FnOvZ)�Y"Y���y<�l�෸~贞�)Lߧn�h ����Ǣ7����b{��"�J�K����h�@N��1�a�(�Ո��n��nmߖ\��N<��pZ�?�F��̛9�3<r���->����2��1GDPo�]�}�{��[z���~Bv�8��uXۚ��#t�
�*��o>�v��f��Coq�ٴ3~��[T{34��$xZ�Y١����V���0��hE[���C��3'�BNl2Ծ{�kX����S^5�֯�os\��9�Wg	l�8Ĝ���<2y��sX���AטR<����O����Hj8��Жiv|0��O�|ɨG�C�k�3U}�h8�O�*�Q��Rjc=��Ԡ�IB�:�����Ҝ�'�6��W���u��IfIߙ�	�p��$��/,�@�+dG����*��2=��R�T?�0��$��'���oѴn�Yk�]/���Bwx�fJ���U=��"T'��gAQ��@���阇���r�_����,-�� �'��g4����/�7�S[/G��Ft!���u+hc�X��T�g�U�U��Vm*=Y#�V�G��m���\.�K3�
���=V�ʌ
AT|�6*�<L~��e%m9Ow_�u��������ś1��v�QQ-~������qޗ%_A\�ֶ۸�'�q�4���nQ�"��S~em%�on�<'�LG���%�ܷ�(?;��R���:Pr#!�E'+���)g�8F��X�R9L`4�-CU�C����2n2*d$҉��c�T���a|? 9
�р֤�*�C����J�I����UZE��R��A{����J�[Agw�C�����lhs�ꐁ�d��}{;��L�t����&K+��ů�,�>U��p�V¾��f��(�F/����K�������O-OD�'�fOa�c7 º�?�m���	o �=���r4��7�0��ZD�'�i�8��8�I�`Zۏ�Ŏ�[v�4��6�� ��(aFӃ��Ra]�U�]>��t�2��i�핢�B'��U����������h,�gQ1'o��B��g�T�E��QxȌ���Z�w���֚#y�4?��C����,���\K�Η8�'�p$��т������E2�\;K��� �_y���S��l�f`BkV�-��#)P��ң��|����0�\D,��(+P3���1��\�[ЫA�����AV{��޻W�ѓޖ�~%?]~O�e��Ɨ�����k�`����Tl\��{d
�d��
�|�Ӎ���p-U�d��9��\����E`2su���!f��;��ʋ�w�ف�X\ �2�"�9��nSp��`SlI���P�	�3��P��kq{j�˚ �h'z%s��oĶr�4bU5��~�1j
gʉ��H�ƍ���:l�r��͑O
���Z�Vam����T2�P�0��.x�e�� U�!GSRϼ�<��%�7J�$@�'�p�ԍ�;�Ʉ�&JP��q=c�gu�2�&�*WQ���%�Ȓ�Uܾ,�N���Ԅ�:�z�˭>����2�4�j��~.��瘅������	������KX�B�^@/o��
D�]�8:Ô� ���7�Ʋc�X��f���U^�k����@�<\}M΅M?`6 $ʔ��7��3a܉�*<wZ~��G)4���e<����U��5��x������&�C1�E�߉|��2��@S$&��#r)�[o��8�ڱ�z��F#�P^��@��h+ϔ}4T�_�t�f���Q.�F��7�O�������Dԕ��`7c��c��}ɽso"��a���@�uo��Y�qJ̱8hK��fJ���e��߯?���|�h�������j�u͑p`�4ݎ���-��}XƦp"��!-@�������N����6�b�:Ą���,��+D~1NP�;Y�.^f����.��<2��>&LJ?B�E��fBJ'����<Y�`=�X��ڕ��c�V����ǆYz�׊�a�E�m�(gb�klQ�4M_�k��`��B5L~����m�z����j��Č�h��}.obt� �<�1������0���6zh�h�w�(f�M�]D`y�-k�K%"��[�@��œ��1�*��A��'<O?d�;�v�i�{�xɑ^+?G�T�:3���*�zu%n�xvU]�NTm[#Ve��z��p�SQ�3��X֑�_Y�n� ��O��M���|J�/ms~������ R\�I���B��(�y�5�W|y�+G�&�QN��OX��r�N�j�8����Q���r6����/^P&���p!�-M;�X���	Lo>���r6�HS<�
�N~���Ъ�d]ڨ�+`�zRX��	���\�H�B.����m�qv�9�b�k���Xv.�
YM}.��.�T���V��u�!�mI<���^RJ#���y����J-��
[Nȍf���p�`���0s�E��?kpKt5H�'Z���1Xz��
�1�DNw�����e�����ܹ{W~��ٛ�Y�Vg �d������&�b�ބMM��IGN7I�j��E����ŕ��"e����`:V4�C �\c]���RC"�R�,J��X��ev��7��;�%��X�҅?�V��"�>.tjK�+��kh��C[���yp��pƸNp�7�e��ϗC��da�������u.K&o&�7~�Fj�gO�(����R�ͽ臼��0hQİʚs�U/+�o}��5}:i?���\W�j�lk��b�]���xS]ג��K��Ë._���T]�G�.]\���[/Hx��U������	x��yÞ�O�;[؍a���MU3�9v)�A�E�X��2hq���f��û�P�A@��9!�4��+:z��rWaG#g�����&60�=�?
l��,��T?�G�Mf��"Z���8I{�AUa�K䐷��Z��=ID�6�F�������d^�S}..�_\�^U��ߞ>m�oz��j@7qZҴ�ʳJ��pU��3����҃�ݐ��y�m��;*���q�ԗ�g�CK����Nє`z	>e��t������w��XL#�2�v��r�(��7�~����(h/����mx��pq�_.�-?�u��(l e�A6����h��57l}&�6jY�CY�3�:-x�<T�;<3�ҎW����M6= z'��
ѐڴ���{�%*m��9E��xqe\���l�`�B��I(�����}��&Qo[�Ƿ��Z������U0��V�ʾ�����3�
nH��:Z�cr�H�o8H�q:��(��-j��T�OE�c��J��)�*�6���@`��:����-A�0v��(�2��D'�w����hzK�}��r��F_V�h,�҈Z�ņ^۝��r�
jWAG�/+�l���)���d��x+$�0��r�H)zyNB�P���l%�+���5����nP�t[����z��d;���J;���A��i��^�p����h�.�l#J\��d��ׄ�\:
S��׎�����|�
��6�uˬ'L-p��y�N����'��@�2NP8݁�d#��;ec�y[;�K����6�	A�ۦ�����x][a@_h��wKC�M��bG�JMk�(�J=�gA���ut�ua¸�ݻC�H`��og�+�!@L����֒;��l�H�A� <1�ܮ#>b��I�-o���=ss��|�5��f�V~$���
U��	8�o�{����N�A�ձ���8e�����F`E�_e�V�/�ג�J��%peAq*B��p�ߡ3c��I�L���K3֛�D������q,K#�u���Q5��� �R�z}X�E̩_�'��Ŧ{��0�LF7�q��o�nx�z�K�����c?��C X���mp��1fi�hx��$#_MJ�|E8�j��6D���Ӵe���# %�I'0s,C8�T�j?c:76�����ٖ،��T�3�v !�:#Z�����W�e�|��?�Wg����|�P�r����q>`�8,�uvN&��Њ��DH���2�ؑ⳨!dЌ����g�����������Wik��@�_5:�o(G;��-�l4K�c��nر�;&����dƒ��.܀G����X��O�16SF&ZJ9J��*ڗS
���84�Rc��ꛤ,Vj��4�)?�4��� ���<���l��R��Cp���e���?����+1�@��u��\���`�v�X�y�|R ���V{ײ�t��H@Y�R8h:g��T��]���n�������2�Ճ#�q�T;i��fKM�0:�D��N�F>s����������k�oU�����c�!e���O���ѷ� �$-4q����lاV �v3�#ѻ
�KA�[���M�&Wpx?'m�$I0<�,�\�ݍ�u��f����m+�7��&�u} s�8��x���e/ɷ��X������VbX��0�0!��1K��/�
��I����}�=�;Ca�@gM�7+����gl+FѯAzwt: ھ��cb�}jZ�۱�Ēr�K[=@����,�ϰFr��T������6
���b��V�j4/�&�昪���4�����&yŤcB~�4/Qw�;�.�
�����W�UE�L�Hg��D�dp��j�Y��w�M:��.}��]��/�/Q�(wW�����֩������گ�����E@xux�N)/�m��Bl8�}QV���B4��n\�K�m��"�d�܂3H�Y���.*��w�]qӚu1|	9lS'�6������de	s)��B�I�X�K�mG�YV�� ���0L�������oKR���SY���Ħ���Zs�Ee���/2�Y����(��ث��@�A@���,�1��%�z
�Q�ʡ��QS�J�+������c���n�P��
`�f��b�]��	g���� �&di&��%�F�C�U���?�\�P���:��\K�L�0젽JZ�Tl/Q��^M�(�L���ʡ-_h�P[��£EE`PZu>�F��M� � 0Z��Nlc_N�c$ao���` �;�4QrBe�um
��u�����й��(�$���
U�E��%=�6�&�(OSVԝ�xN�J���F,TǻC��g�	J���~�S����{�D���^5@V��U������&�I(.ǩu�.�*}ǯ��ԑ�i<�}Gl"L'_F����u%�\��u�S��d�WY[��/�ؙsi�.|����6QE��.�Z�����y[�R�*�Fd%c����ۦ���)B
��Z�8+D]�����h�(�#��O��#���sρ�S������ః�m1��&N�hK�����;����`iYўl
_Bv|��C1n�_�?�E�'{&h��1��Y��.4�~MG��ĩb��R�2'�.K�oy�a|�Ϧk�ژ�V���N͊��
�W��Wd=N�@p���w���m�s/1�^O�)�Ul��p<Cd��B��Cc5f��^*�Zr����P���c�y�ml	�RC� ?Q��K��Y*
���5��<��Jނs�%<�(s�����N�4�DVU-z*������z���м�l	r#�m�!�>F�ރF�Ζ��;�� r�|n������`�:��P��Y�2�tM��/�n������Qsf9T��޷U�WL������cY rW��)v��#*h������ܥ�&p_�GT
�ۖ�>�.��`We�&<收3
o�'��lv��� 	 kꉻ�B��rGJ�b���_�ƴ"	��`�o�Mݳj�N�q=|�W1�ts[^�j���2�Z��\W�R��W�M>�O.*��}F���{�!!0U���t����h�O=Ơ�Y���:U�5͢l��>/����<��x#Ɣ;3��0[�w�΁�b�n���i�	0/�W"�^�`����_f�u�����ci�E��U� r��D�����C3��qӡ��9u��H�2G�1
��KM�d�[�n�7������1=���������|['B��2�&t���K����p� �����a$PO���ԇ%|m�Fa�.*q�%�%��tU���?�mF�Z5&ɔ��4f-k:�Pn�,~��&qݛ;����*�e�����ht*g�fiY^&{j  &&��A@��j$�%q<�V��Ff���%U�OVK�����I�����%Dv�c�wq`�_M�N��d����	�>�{�ôV�[aGM���~�2�j�`%��g(0,u�m��}�P���b���p��|�3��;�b�mM�ke���~�ƣ7��@�Mv�ZSԿ'�Z;	��r�0g��9�b���c�h��YRHrj�Cw�W0|�+y�x��u��a��I
���bk"v�F�4�#y�]1�=6Ym��	cJ18��f5�)uN[Ŷ��_`l��_Ts��C��2'�x��I�_�ҖGy%����4�}k���!<�tF�=�]w� G�Fk�ۭ�Z�f�#�s��Ւ�H�%QZTȉf��$�I���x+Tk��!�A:��{��muop�����#}?�&�����e��O�79��M8X���Ʈެl��:E��sp#��C�<|d��N�:�c�cG���U	�O�]'�VD�u��<ѧ��M޼���ͩH�c&��<��� Mjw���Or����
�~��#}S�w�g�֕�^84�Z}�~�îm��@�Jk
��^^�L>�sf�?��қ��M��Yb.�$֓�$�#���y?��d��h���PC	����Pg�e�G1$�/
B�E,�����`ke,���wMX�I�0Y��/�7�qE ~���l��yS�+$mϕO�
����ϒ!�N�m�QS�:��O��'M�����v��:���h
0� �ݬ��L��\6��K
��K�	»��=+�ܿp^�fK��=9��������W��ȗ�N��+�)�$��˓-�ș�2WV�
8�v�[�?b�c���0kf�8�x=�5bC��3��Z�/�B�x�]��	W�JV��k<�r��9�Y�~T�{^w�~8N��Ј#f�� =�P�P^�3�x�o�+������[�;�'M����d�M%w�;��S���Z]	Ř��p�<��	�_薥b�� @�"��M�K���Z��aQ�P�sF�^D�eMI��Yyd�8mEL�r�1�=�l�x�ڛ��#�	�m�b�w�P=ѱԢ���Cn,�8��9k�=&{̦z$X.i��N�\�|�Ȭ���y��4�sr��v�@^� K��Q0nǪ���y���2�+	tM����%"&B�`Y�_��I} �lְ�Uiۛ���H�n{�yL7Q+��˸���i�λ�c���8[�KU��d��C�+(R6ݝT>M�0ՠ�kp��ԸM�b���*R��19��O�k)?�!�U׋'Q�G���P��ʂ͜�~�
BR���U[�m5�;��n R��9�9��������r|��3�����S�|ý�DRA��s������7>%�H����K�	��~���j�nԧ�M�2�d�G֏�FF�t�Z�!`+`�'E���\�#�NY���'��1���ّ38��� �wf�tv��<M���,�^��%�ؒ�+�������s�Wh�˯�2�P��إ,/�Rs?���]�\<̖�9YỿK��[W��!rtUi�"F���9�b~��5�󊦎J]!�mo����
�O��ݶm��K,#S��*�
_��=k_i9�O ��"�{� CVq� ���mT>e,�� ����kg��[��[;�H�(r1�']er���G]wD�|�&�z^�қ곭|!:f(S�*�80D��(u����x��h�t�1v7��$ E_�s��w�%W��Dx<@T���y�V2�D�Q��t&a��Щ�y(���F�T��쉪�tΥEj�
t��Xr�S
B.��(�T�L~�© �!��uӫ2@3{�
g��hB8�$F���G4q��*��7�;�G"�z�U�A��T��RWiC�v��E�#E	%������h8�c�ݡ����Μ,@�j��j��/�%D_)����j��ʙB�d/\FT��4)��e��i����{W&��`��=�4G��~�t�K��9�1{6!,_8V��we�k��ʠ�P�:���.��Btkѱ�:H�H���I����Y�c�ҟo'��`������6�[Z�j
h��l�J�h#9;B^;/��TBA�)��k��s�Ր�Ze��Έ�d]:Km�xu�G٪��t6a�����E	��=�����#Ǽ�m���Ny��#f�Ɣq�b�\�T�����V��G��7� #� �?��;WЯ0��pN4�Zo#�!/ H }{��R�u6�vE߯������B���il-��D�)�s&��z��%���k�"tЇ8	tj��������9Cpo����Γ��c�/�h���ҏ08��Wzj^5�0a+h��5'z;aJ�8�P���KuJ�����X��]�p��$�j[;j�������� �z��ia�O~���d����;�w}"(�H�]���"\�u��ǩQ�i$��ϛ�8�%� ��lz#����hێO�w\��K!5�=n���&��!v4���LЕ�0����LZ�z���ܥ�Y�{��K}�5B����Q�d|��
ܚ�G�U�p��� 6P�y/�+���
�&#�K�t%�<������Y��#��k�! Bb���ذ�d(�!���*E��	5B�ϲ����ʷ��[��<W��N��7���5���y�m����r9��џ���
��H72�LZw���4�|��S�6��8��;���1k/�/I}��p���N�l�e�'��^N��;z{��q��)Y}��>��N��nh�Զ8�����F�t��2��]�>ν�<���^M����D�~_ϐm�?���ؾ���C�z_Rn��G���ג��kz��h�[��n��ݿ��@+Mk�������4L6�{J2�8��+HUO�����>_>@{@E��M�Y��/'��u��y1Uz��i���3�Q���t��ā3��]��0��-���7��>��)��>K�p�������������w5[{K��S$�`�.�y{	�t�n��F��j�W:%���q�>��X�-�'�g�Z�� ���QgB]����mS.90�
Mu.�Hcs��t`M��S������V����K���-��.�7�!_�2쮤 ��uϴ���v~a�O&�N<J�X�1�;�E*�\���)����e^%OH��R�}����k8w����jx��}�cJ��]5�gܥ�ήٵ}�*lDm�^��D���}+r����>�0�V|r�:���o�����~ϻ�{!f#J�? �B���8`�x�ȱc���-ӹb��E���UQ�QzC�ҕ��-��@ �n>aE�ϥIe�y�X�R�'aZ�Z4�`�
���(J'����1��.��h讇�9�qZ)I7�l�bz���Mj�z��"JQ֬�W}o�̘4���^>�)^=��]8G?��m̌�՟pH��*�i;�fEcWZ��	����j���u�"����eR�*��a2X�MT]�P����=Gly���_�b<:U�M��*�,{$���i ����7�χ�밌��p�|o�t^Е8����[K�bP�/PV��|�	I-M~�ʬ�qj}{�8l�%	�&��{o�I��O��l��`"}��~.h\f#fL�p�:4�D���I.�1�d�ҟk��nyO�K���Į4�G���:&�ٷ�$E�y�g��
�S�ux���_V��&
�fVA�>-	.-ioo��'c��ۀ�Pr�;���$��duix>�8&�o_�8)�+�y'���[PIf7��?^�����R�ђ�5��]�w��@&��#yZ�2���W5O�z���+J:U��DD�3�R�0:��lԷ>x67�M�1B��NA�OKT����1�J��DR�����L�ɑ�P��k:qWPПx����ś_ߪ��m�S㰨��4�ӌ�NX����Up�O�
`���S�ǖ����7 ��2�wV���wC�#@ � �ۃYM�g���_�`���Γ�[C£C,���2B�j�SNcc��>�i�Ko�����c�l�|��N0E'��ioTsq�"]�!O�l�5e��[C_�P�m��b�$h����I�g\��8V߶�,^��#TkV�E�g!'GΜ�3/�&Vc6��<� 
MG*Zh����٪>�L��q^1+���j�$P�J�l����vS��f�N	�o����AΘ"����Π�\��IW�����al,m�M]q��g�.6��v*����
y�"�Fѵc�D�!˲�u{���"8���x�J96����p��DW��w�h|�ȶ5I�3r�uڙ�������v��NА�oS������ڈS.lU~]V3���K�6o�m�$m��9R�v��g�i���_5��2O"�d��]Y�Ȫ)H1k�`o9,��/�m	i��5�im�|=������1'&��j��7EKC�"S����q>����Bzq��b�s-�
��b�á'[���s�,ś�i��#�xZ���%�;�y�p�cJ�{#='B��L=���+z!�±_>�b�G�M�j� 1H�B9���ZRxn9, ��ۍ_4�K�g'T����Fkl���a�ږ�?�H�/�0D�r4,O�G�c��r�g��;÷�@�5���x|��e2��Tr2�-x��5��\�����/�dj��V�� Sוi�u�d!Q���g�O`����(�F�x��=;�Z�cg�ih����/�f���mil+ږ�V�������������e�,���+��ů>��H�����?Ř����ۢ�@�^�����u;�����[>�/,��&�	������^����\R,6{�5��Y~��� ���D�ٛM�Ͳ�Q��w@�-�z��dV�T�|��4V�U�K���a���gm�"��ȇ��.�P[Fd���⮚���ğ��z�6�[eL�п}S�4�n�MQ��r�N֯�xi��INq����4��H��CG�$S�r�2F�]3�<��h��q{�|p��[����>�F.���*:�	T�$� ��ۿ�'@1����H��\)Ϭ�
5z}]��m��p��-�����wh�7�ȵꝦ���f�ѯG��4�h�}^�I���vP�HZ8���X���b���w�t�X�A���b���xXE����~�3
۴��t�ePgR|�f�RT�F,�ؐ�{�@O�vl��l@X\�q��d�����P�4�C�!��)�5��u޶s����$3_�%$>/����U��l�|���/wk[.`�/n�qaKy؝C`����1�:�]��I.�e1A���N"`6���X�Bd4�a,��/݀\W��X��_�L���װc2�\X ���bFi� ��_����u;���Ɗ| 	�)E8x�N����]D�޿&9��*�u��~���SL�x�˭2О39��"�2Es֓H���2W:�̍+��J���؟*	�Z�v[�@�G��T�/��+�5�K�����Tυ��z�jA�����K�a�.��ȯ�,���Dk
��2����.�0��{B�ꆽ�I�30���5�r�\��ѿ��:�F�[ǵ�c��@��Nɡl�����j1DS_}[Kw�Y/y��s4k����f���C�_~�ٹ���?���G/7E���GdF3l�_ Ը�,��?����s��޻NW�m�r���DX���_uJږX�8��3��7�D�#����_�7`�v�� ��D���9��ڃ��[!�Do��&���x��(�g���/�r�a�Y��<���Q����Cx��}
�����q�J��"�<��2C���?�x�$��<2���6h-
�N�盥)�O�+�7!	�XT1.�9��n�if�����a�T�qa��v�Z��3��6Y$tB��=�S�[4;T�Mܦ�X���q���)����%��U�ݛ0g����-*2C#;3��?��Κ����ŧ���#�׷UkMi��P?�>s���͋�-c9�.I&�B1��S��偵�ר~R�APWa��m{��`�r\��o�.6	1)�Q��DE��C2b;6Z�;���%L�K0�����3E���+z���̧���[	/����F�F�t�|���U��;�H�.>p4�vo#�0𺆙QruikfʏW�%�C����Y�]X|��w_"�Ŷ������3i/�"�|c���Tm��_�B��L�Z��6�P�%>a������k\��ke��)$��G=���Ğ�#�`	q7C@�b�x����G
������>�V;�}��2�$�OL0I��h��e���R&���\f��A�jo��m��pMaD'�D �qC?����0#�l�I�n���%R:�jJ�x���%?���а����b��tG_��M4�2������_����-S2꽆�0�G��L~�b���� Kf�rSx�U�SWҗJ��U�&$�{ ���TIu��ǵ�c���c+��nyF��(A�U��Ǉ:�Qg�|���+T�Q�X|Ŵh���]I��A�h�(��?�7G\Ԅhl�!L�y�~����Jw��IH�a��ū�8건�����	e�?n���x�>��C#���ѧ��s�CX�5�t��/�2S{Y9�2'�L�j��W�w�!��'$S��d���M2�4,4LA��)�į�%i���Y��b>A����+�d<��E!�d��I�����6!�-:7��F��!&�h\�������gQz���k0�%��l�$/&�vaq�ME/l	�І�Eg��O6`��g�?$�7+ީ�Xi��<	�]I��*+ &6J��˂��W+�4��%H�f5p���J�஽k�����2Z���C.A�"�Bl
lRa��OA&3s�$���]�Q�~��1��F�n��F�����M~���bn+���VN�p~}���}��[�ˠ��-�%��ڵ}X��K�O�ET�O>u�SN۞�������CD�������ipĖ��������^,.���k�����rߍ�`���G&��m�aN�\��'L1�E�z�9Z[�dW�~oOV���Gn���x�r���h�+�e
z��T}jݦyuMSK�8ץw/H@I��4�B6#�~d��t(�����2Xn�V�>,���[9Js��/
K��-@�F��;�2�;{"�ߝ�?o��%h_j~���͇[n�*��a�)w*��e1ȷQ#}�����M�n���k^����u�NW�%
@/��a����Cs��4w8����15A"�y�BM��1UG5t &c�"��콏<`ǈ+�m� �W��$�N���jZ��+� =`(�TRH �L$�g&���=�5z�2�糰���S��P̦t��+��&�h�f�s�Q}��h��7����D�/k�voVN�xT�Z��vؚ����s��S�ۺ�A(W0���sZӌ�����8�̆���S�_�Tˀ�I\�� �zd9t_�p���n�hj�^^Zyh���uo, �)��	���a�(�X@��f��-j'��Ƨ��0�)+�=��X�#��R�d�g\��PҁU��C���ׅ�<����Y<|�\J'���ig��΂A�02y�B>_K0�ӶO B�N��,�Tf�=x�{v]�\�v���e��w���S$+Mr]S�ixs^��ʆ�S_�x�0�������I�u/~�K94�K�d��nA�m[�i-	�n�<�'�Ƹ4A�"# �����1̈P_�s�B�`�BN���%���$K/h�=���X�t|zd���
1�`N=!�N6�#��/�����N������7t͕��{i֎��#�d}��w��7$�w�+�����+bxĽ,!΄�А�]��8�9]��Mp_;����^�۱s~]~~��DU�S_��q�����?!���beU��X4�)�/Ӡ�6T����{o����xk�*S��)���O��/�����A>R=�Ԛ�-���_v�S`�k��w����U�ol�w� ��eD�&B�s�w�y6��&��^���.Y��VL�W�����m��Y-%���)��]�:[H]N!�қ$�@�"���Pg�
Z��Lb�m��TUqI�XZ�0/���Em�oQ?��ƿ�*������'hP�N�|Q��W�8�7*��@Z�!��"$�f�=�EU~Ζ�l��e�6��xH�o�w�d?,P)P��������m��~M����z�,)K&*�{�� G�hL_%?� qB�
���Tܲ�8���)d:
B�q��`+�F����������5Z��)4���@}�0�iX���.E�]p��<&�T�7=^�bP����!�] �]�>�;��P��́��G�fj�D/{;|	��yLb'�28�T��lؾn�]R�b\V@[B�c|H�u�^[���ƕk.~�G�vO��si��3��$�	^�9/�.�B�z���PF�/�U���qp|�p����� l��r�]Q1覂��#�L)}���c���� P�W��p�������⦑��Q���֏��b�{-�͜%�-�c#�N�љ��h���2��z�.��=���>��ʰ�V�)��գG��^�XE&v^��$8^?�_|'�E}_�%�C0����k�am[�U�Dz-�wӶ�b>ͳ�9��]�����h�k�mFJpH[��N���ǦO���ߎ��S���ap	�k�<���>;L#E�D�qy����=:��JRM4WO ���q����	q>�?�e[m�8�0���/Y�L[U]y���|����s3�����B9�4X�)�>rK���4mS��G ��s�ݶ�"��Q\��w�8���x�}iXt��0��#�'s[�+�c���,UrM�܅��Y��*�$apjjh���5�\��2M��|�@�'��j�	�N�p�&�B�;�<ܪ���,Ȧ��P'5a�Y�m+�{�G����C8�d�x	�ޥ)�9^_�pGR8�\�aO�ّ�s�����%"���],BKׄ܀�@����ʲ��}ݶ�m%�kۓuwU0lh�^�iAD_پT�����o����T�i$�*�Z��у4�y��(�v�W���1�p�R����(ݒ��u��P�˖�V<k�%QU���X�����]��l�V0�.�0�t��%L�C �8in+�`��H3��b�leo�7.b�]gC	gU�w�9��0Ճ��s��a����O�^�f'�ļe�;%�g^rS��Y��W!5ެ��[{��~�\j5Ov�������:
����͓&@7�xշ����a7s�:/�(:�P秷��A
u2��ܕr���wz�(\�{T?������"������7d^���ȇi���'�ݠy*�
��(t�e�Z�"�?U�bj�i �:��X\u���I3�����d��骝`����"���(2N�Mv_�O�������
����_!*>B�b��3���&��|<*�a6��,$ᇠ�?� �#yj�a��Ժ�x|��Ȃ.�Я��0xEe_��s�_�S��2`��C�](��Dx���U��כ3�Ȓ��}Vԯ�0���_&��=�����Z|v!-���?��썬�/��4�4^�W���m���|�хMm3��c�Lю���(`�0�>�8�Ix����P���#��+�KPnM��cH�O]5�K��7⢁��ഀN1/D �ӳ<�pRAy�lf��>\4��wK� T
)�x�o#nY6Tfwf�3W0HP
��:\��M4���7a�S�/�#���A�� � �>��YSiR�Pd�cg���Z�mi��~$���G�f"@6�x��	p�e����J���r�D��1s4S!UMu�,��8�n��f}/'߁������+�	�'�R��[��!�H��aھ�^(�<tջ`�$y�o�8�n�a�?1E��c���%bj>��bD�q�V���PP��)��S��b�E�� \G�f��2�$��W��Qr�(��v�Ɏ������?g�K�Z�,�3.�f���
�?n\;���:z*��bU׌Q�\dR}@�L�m�!�sV���;+�ބWFY�*�)�VJO�zTB��}��u�����ʑƒ�6_0e��5��2Buy�J���Fn�I�G�k��p��I�N&B�а,҇��y �*n֑7na�zf���rɩx_#��ɚ/l�0Ӂt��(dlK$Z�xi�Z����߲�����>�ak�����Ժ�{%7�������A!kIɺ��((�Ui�
\�Ɛ�QI�����a �eϕuF����0�F$K�����I�jj!��f���L[um�QZ�fK�l�`�AL@Ho�G��n�+L=I,���IO��&L��a|�B׬��Q�$��Rap*ܕ����6��&�Om�C/�R�D�
�(�Y�ޞ����r}���U�}p�Q1LCx�_�)_W����i�e�zG3]{������q֫��2�������=�%Y2�n�	G|DE�v��9�����A�*��R1������ڿgC��0�𦦨}��ܞ���#��֮\F�����^%�a��s�Wf���˫�q�y�k��U@�&)�6F��'®��I�v=!z���/����ߠL[6;��W���X,rE3����i:����l��	�� +�+��Y�� ������VKs߁2	0��C;�7)k�N�ɏ'u�K���( ���%��X���O�XC��{�ٷ]��t�	���ȯ%^!�+�S�4��덲�5�M�c�Р�"��T��|`i]��z���ip��@;3ڮ��h_��0C�"����~h�Vk���/8"�w�l?�������0�'�4Iw�wLawd�!a� �ԗGIOՅJ�Jp�ɳ�����h�ؗ�>ePȭ�ѪNm�,ׁ�}<U�:\@�kJy����"�6�*!�N��3�E<t|:�����n,�x�^ImXX�����?F����KM^H����H%�s�P�n�oE�x��O=�c���Y��7u�MKh��[�,��/B�y�y��奿�11�h�>2U��
֞i��V��w�,u�)�-� �RrޘZzD7��CE�	��r�����V���|������F��3�i�53����:����B��-�i$�@�l�pMv���1N�j�)��u���*���KO"���z ��E=y�X>�[3�9���`3ږ����kS�;���TEc}���f$P}ٞ�ie��d��d�(V$�a�0u���������د��x�%�5x���j��B�jbG�(�5��&2��Cx����;�i�~�j�o���Ӣ�`qh��u&��K���Ep��lI�G`y�8�(�K϶wV���ߪjFx,`�ZO�ʂ�&\�y%���e�W ��ǛG��Dnp�����nM�S�����3ܻ���	���L�*�-���+Z�c�P+S˳�|����|���V-���c;i��Pi$;��z��QMw��}��ha'c'h[I���:�����Z���!/ɉ�>M�xV[v�����}]BPl���_��u�p���e��"�c�"_�7hY�-A��洛Z�4I���?4�ǭ�M�n�r�ǣ���I��fk���x����E��&d2c]�:�=�A�4�����g̝OSo��#����x�8��bp�=� ����{��f�&�;�ߴ.��K=J�/��^|.m�F�1�f�B��4�D��?�&RS�_E�,VFʰ�|å� �K��8xyK�tS�B�Y&��h��Ff<��&˰�X�9��`И�+?}])���H��蛂�?h�B��:e�8��<�����¸��u���ʐ@Pz���� ����cYJWv7]0��;X�N�ǡ�C�Υ��k�̙KD/<x�<�K
l�J$�~����sG�<��W�ժ.�Q# :���*�6A]�Q����{z�}�!�w��!뛍!
x5ߡ�X�]@l��fN;�����}�u�G�fr�!�4�0_���R0�W�����~�H��r�D��w�R&��`��9 �lb�7���e&Q�ia(�M�^���U�τ٣��I� ���IZ�H���V�w�������_@��ҿP�Ch{Ie�7q35=�����(M��
�`l���}5�{m.�������(���`��\�oF#�nA��T��M����s�-��>���3T:���$���(����l�q����[���p�[��fG�	��(?�Q|*Ķy��?1�f�Z!��
��]�a���v"���c�4��u�]�1u��|Yi�����=�~�O�C�k��#dМ���n�!'��d{j0G�4�v�ďr'rF��Yy�A;W��<�>�TI�/7��K?l��`�/Pm�ر:�5�5������fPaitО�%<W� �+F���U���: Y��塷<��H�����H>_<u1�t3�-�{��4��O�HK��g��D{��\����8p����6n<iHť�r�K,�B嵡!7ۂ��-�%������O~Af�3rp�︣ș0z��=w�0w�1�����̫�KrE�T�j���w��B~kp�A�<F|Qقπu��(KUyq;�H4�w˺� Y�_�X��c�d��	��1��l^�޽�e�f']�3��$ @<�F��N�	�R���k��Wy�|~&G�6=�p-t�߿�&����ڠ��Ɣx�|�\���쟍l�����!�-������\��J�9M�>��O9�ۉܢ�A"e�ۗ7s�HY|���(�����Wi�y�ve.z�Sr�����^{.>T6Ӭ�Ț���A�CqЬ�hP	,�~�jqFtw�5���k���`h���L��i
���t�x�^W,�a�n�v�7��(����jKN�~ɟ��anA�U�խo�nq,ȅ��M��tb<�z��눀/���;�(r�=,����-}Pk�:ꪉF�Մ��(����� �j��-o�c3כޟ:A䖁}X��L�kOQ5>�*xj)C�R��4%�5¼0�2��Z�Ӎ�N���"J���Y՘����zA�$��-,#���e���dʡ�P�}FrW&�Q��J�����M�*_�F̜��ѵf3����Tfc��G}q+�[g�D�o��UC.(�~Y ������6Q|8�}�k�#���m>��`���0`�͟*�XHb%�xcЄ��p�q���u�|����#��l8�3Q�l��3��‧H�~S���Y���6u��Y���O�"��܎�R�<S��\b��t{RGqRtH�b�k�׋�Aqr~e������@[G"{:}���r�{_.�Qhr1����^�UPKp�"P'ঃG��1 !�g�p��Om�������*W/�JEz�6J�T,���8����E��嶙�Y�X��8I���o���nY����^H��*x����P� ��T� j��eN�3��*w.�_�ᱽXz����+�vI���pX�UBv�̔���bTEc9i1GxV�'�S��	��yV_�+����\؈{�j�@�W�n�@���I��.�7�P4a����p�i#�#��"�r��z������ �C��ߤ���Q͇�����ƹ�9�?x[�Μ��q��t��O�l:<H��x;����S	_�6u�! �9!yIm:W�����	�%�M�,/���HK�7�#C��29m9�	���k"��2���~����5�ӻ�{,����`V(��cC�k�D����{&�2�g�6�J$$s"D�<�����V6�)���21�/��xj�ܰ��{�
D��O�<H�A�x8���V��6M��ǰA��k2�Uh1���G6���ȩ���l�u���
(�'�9=�xv *��l�>��U�����'\
�_n? eQ��^X.>5ŵ�fb��� :"����89��e��hQ����K/�c|"�]o�˝D���Ci,A�u>v�*��*ϋ$�i8�Q�@�Vt?�H�ѹ�s�"���czF�?Sb��v����%Q��7\�:�����P����=��kP^I�^N�נּ�6z��Y�� Lm�ϿhsL���y:e�5K�*=��͗��3L��� �Fĩ�'dvd��jb�-����.}:,��v�t��geH�T����R�J�}��'���Z� iĒc�K�����`���M��ʗ]`ə���[�"��W���B���·l�a�{�����O��,MM��QT�A�*'Q�ɧ�q᤽8��r�x����v�>�V�����[�ǋ�����h^���j�#�;�M�OR������"x�H㹷4���f��G�zB^ ���Q ��iј�1yi&��wT��B�h@� .4Դ4�<�6O>������H���f��
���w#!�����X��:�Lj4�b���)7�l���s�d�5�wa%kp�dݲs��U�@�B����ٰO�#�c��v��z�pm���3L���e$ΰ�5y�-I�d�LsP�J�/H�uˁt5�?�k���������̢<f�Y1�,Eq$1�1	Y���7^v	8�ΰ�� !����4~Q��Ǔc��/{I0m�g��#�X�H:�ΰ4Z�g�'ɺz6:J��Z�`t�c���t���;b����W\^�`.� V�:L��l�cQ_Y��O�K�ls6��3S��}c��]�,��(J�ޥ �'/������lZ˫���nӂ�g���J��)+U�l�E�eB���+OP
��zc_j��GDS�>2)|�5m���	M���k�WuE�E�!�  ]�x��X<0,Z�g#(<��,�掁�{�����p�E���t�Ja�G�7�ݔ"ܼ��`��&��%B4��|q�_c�ѽ�ʂ�Nx��J�*����@��U�nG_�!�0��J�2G�P��Ҍ��;�J���T��
63݀�!����� ,��,����I��9����e���R"ur����Xf�XB��A�/G�+������M��*�%K0T(q��0��m���B��qͫ�]�%��A>�\��U��=���;5�A��O��ŤJ��z��U$�è��jr]��?O���Gt�O�}��=<&(9�w�f8��A\@�_8V]>c߇:��t���&c� m�v���1RGL�UD��!�2�z�uc����ܷ�����ݨ|�4�����?�J�:�3^�������å�:a������8Ӊ�R��KM<Y�(ڐ`Wa�W�
ۃ~��v ��͙�+m�XZ5�����&�^Z�Y�_�lC�lÚ�f1���)��ǣ�@�	||��m���z�_��֓"�bťj9�tE=\Nb��B-G��A�
��E~
������i)�5� �>8��2�g���x|�ʝ���2��pG�*��EvXsK���X͎�Q*\�M�S"�
�t���'��w�
���������f�~�2I0�Q	�r�g�q���{1�mS+rd�q�3r��}�WG� �JgF���sM9��ńDĞO���rt4��c1���A`%�*�8�ݷ���ş=����Z�=ۂ�#�ă�N]h^�\ސ�i�Ow��=�p<M(|�]a�aA��.	�'d}�����j~��I� �bմ�@H1y��wl�ɝ{�_Ċ�~��V��i[,�K�Q����Vr]��0��:��I�3C�7��M�r�C�$�/({�s�qٞ���|�W��r����]�A#�(g��q�̤R�|�į�����}�Dї�7�tMb�8�"��G�b��0F�E�qO���?@��lx4�̅ä�)��PJo����F��l� ������O�N�M�/� ^],J��=V4V�%B^����.2�U�R7F�liz7p�Ǉ�Od,�x*����j��0�۶"��=v���c�t�n�}I1�r��w퀃���U�'��M��9�[�)��H��)D�uK��s�n�&��T�?#���� ]��������'uh�?��^>���>q�F�Ky��ہ��0�����F}֥���`Cv��n�y�β$�R�yt3���Y����WbZ�w� �$_���eR 6�|�3�������o5��g��v�T�.�<*�.iO�~<�=�[�e�1���oI�R��#��j�Z�?w�b�}��u��ʸ,��$�,�<M�teʆ\�9��Y�Yy%Xqm�|Gq��J��-���~�"��U!Er��ǈ�BN�+����u�$ᆀ�d��W�T��%5RA�����!�x{�X�V�C��_R`Q���tU"���TQgA����h51W^f'�)�;�J �d�(�g�ڝVC_:� ��6��$��7�����9|�A+��5����@C]",%C�%��J��)2-��.����#ŭ?Rӱ�'�~���&^h�qt��{��u0DF��!�ٷ��4^���o�ck8#4����ww�V���<M����[Qb�iHG�~hE�p��k�{$C�����!��m{�/J��5�YX���u������9X�������������cn��'@T���ۛd�����(f�=nQ��w��Zv�Yu2�'2�,�ȗ��0��7�^�3cĝ�r�q5��vqfJ��(��{y0�v������4"9Է�b��~��+�C�~��6]���qw����}I���QSv�d@��j=�rDp)v`�����qw��SX��(�S��2��G���c���h;�&k(���C���m�[��V�o嵴��.pO�{č]ok�ҭ ����c�:��i�x>]�jh���|�rYc�pR��<*��������i�};�^~ݟX!OD*@+���p���p��ұi��݁U��y��'�3 ��)����hn#�����ں�E�����I3�E���9���$�R�����:nd�����`���_�H�9~�nYI�R�44��2ޜHX>]3KvDe�����C� �J"K��|>���h04����cĀ��n������ �Rx��`�-��[C��Ѩt[����(�
�B�R��߯Zm�Iɯ���FE�p������':($� e�K��`&��Ѝ�X8��F9:NȠ	��&w�}m(U�r�t����X;N���T���@$F����)�լ��x�x�j�i���Z|��U7 ���f�����4{��uw��	e�雂�Q�l�[�C�P�/���7�q��:4|I��_#b_�vA=�d>o+,�8V-vG/x�M��I�<:�7u�Z�z{Q�-\0ì����#HO��T4��wk78�~a$4	k�Ħ� U`sZ)��Nz��أı)"Ϋ��J�U	�aܬ�
B�Υ�!B��E��';̧��)�C�7S�-m8����2_ָ�4�B[�z���T�7��n9�J|�P0F����Wگ�e����~����)_$$�Td���L�#U�a�����/G���n���*{��ɻ�q�b�ګ�Na$
�k���iO8م9��N�#���&K�ד��̧i�ɍQc[���=S·�E=���'�7�	���D��9�����wP���1��^�l��7�IVX��F�"m��^'���#�Pe��>{�����o �{��1��f�s+p�[:�_��{�x�9X��}�q��	ሕ�6�vC�l�3����#����*� 	Sǹ��d`��qo�й˽ml��[����j�x�ly,"�MS@� 	�m�;?���(i���h�f��h���:كK"7�f`�k�{�#�,H�`����X[hpoA�F��D�MԊ��T۔�����z�z2�{%:�����D�r���Dc#ǞO�4��4���m�B��Oy��Tv� ̣��L�q�����3������޶�.�ĺܿ������T��C8�#���SJr	�~]�^���u�0�������*��s���@����i�A�=kM[���)���<=��i�j6Ӣ�a���l�ge<�q��[��vyM�D���w	v�k�ǃ��q��{"��<ͣ�7�ǲ�p�<,LEac���1e��*�y����k�X�i|�u����c	�����v��W��H�q�La�.cݎ����eo�V�V������j����{~��t����,3a�TT��iHu�����M��#�#{`��]��h��t�ذ�2����_�;�,�V�9���{+;�������To�N�$bI�ߏ+l������=���\��0q��8	[�Rs��H��t��;2!�Q����v��
&�@�8� �c��P�u]���p���.��4{��w��~,��_$��T���Ź
���(>ov����$�4&/�R�o���d�R.:Qy��c���Bj����P%��&>M�����h���+<�U��4u�_՞�p��Qj�@�J2�(�-��=���`3���2c5"�E�����kQm	y�� *�R���?4�# ��po��q��'@�w	�3"��af���������	0���3X��l��� =�q#&��8|�
F	�q"�vl�ᎄ�?���øS����m���,18%p>�{*���s�d��,�T��!�Ζ���ȥ)QݹZn2NN,P��]=�ګ��-2u~����KE#\����^習������Qҍ���I�-������m�5���)x6	d���=gd��mfKx��G��oV��Z?���3����;��G���{'ѿ���e��ht�l<�!�Y�V���*�-������-5�ϲ���~X������;4��?�#��^���p5rGt�����i�}x�i�;��|%��u�n�N��-�IH�}:`1N%Õ���T}B?�Z�ﮇj���
��Io�gX����;��G|�,A>FL�=�O� =m�#����=/:p��+�^ܒV��J�fM[�&g�_�C�ϨA������Xh�	n_�������l��a��etc�����:T���������r#P�y���i�lֵ\1� �Y�j[CS��ٙ$MZ�W�OrI�g�e���آ�����&L:��E7�tK'�.��䮔O���3������"�s�Y�=Te˚�p��n�	|x3ǈ{�W��!&N1�ѷyR���
/C�E�oU&^�:~5RV�CP��d�i�P{�D�i�αA!�o���M���"߮�U�:JwT�T=nS�OˌrJ�q�7�(�Ê�Ċ��Z��o:��x4������&��8�i`�Ve�tKEGԾ ,d$�&�TYM���f��)js���~�F&I�ҖB�6�ħm��������� ��yMܺ�ۗ[����WXq��\i�J~�%�Aθ�,7�L5�7V��qz��I�|"